<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-15.1003,-3.72985,138.718,-83.0615</PageViewport>
<gate>
<ID>5</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>306.5,-207</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>12 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>5 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_REGISTER4</type>
<position>298,-190</position>
<output>
<ID>OUT_0</ID>6 </output>
<output>
<ID>OUT_1</ID>12 </output>
<output>
<ID>OUT_2</ID>7 </output>
<output>
<ID>OUT_3</ID>5 </output>
<input>
<ID>clear</ID>20 </input>
<input>
<ID>clock</ID>62 </input>
<input>
<ID>count_enable</ID>62 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_AND2</type>
<position>299,-197.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>296,-207</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>24 </input>
<input>
<ID>IN_2</ID>23 </input>
<input>
<ID>IN_3</ID>21 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_REGISTER4</type>
<position>287.5,-190</position>
<output>
<ID>OUT_0</ID>22 </output>
<output>
<ID>OUT_1</ID>24 </output>
<output>
<ID>OUT_2</ID>23 </output>
<output>
<ID>OUT_3</ID>21 </output>
<input>
<ID>clear</ID>25 </input>
<input>
<ID>clock</ID>20 </input>
<input>
<ID>count_enable</ID>20 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_AND2</type>
<position>288.5,-197.5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>285.5,-207</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>44 </input>
<input>
<ID>IN_2</ID>39 </input>
<input>
<ID>IN_3</ID>33 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_REGISTER4</type>
<position>277,-190</position>
<output>
<ID>OUT_0</ID>38 </output>
<output>
<ID>OUT_1</ID>44 </output>
<output>
<ID>OUT_2</ID>39 </output>
<output>
<ID>OUT_3</ID>33 </output>
<input>
<ID>clear</ID>56 </input>
<input>
<ID>clock</ID>25 </input>
<input>
<ID>count_enable</ID>25 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_AND2</type>
<position>278,-197.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>35</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>275,-207</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>55 </input>
<input>
<ID>IN_2</ID>54 </input>
<input>
<ID>IN_3</ID>52 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>36</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>306.5,-180.5</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>67 </input>
<input>
<ID>IN_2</ID>66 </input>
<input>
<ID>IN_3</ID>64 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_REGISTER4</type>
<position>298,-163.5</position>
<output>
<ID>OUT_0</ID>65 </output>
<output>
<ID>OUT_1</ID>67 </output>
<output>
<ID>OUT_2</ID>66 </output>
<output>
<ID>OUT_3</ID>64 </output>
<input>
<ID>clear</ID>68 </input>
<input>
<ID>clock</ID>90 </input>
<input>
<ID>count_enable</ID>90 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND2</type>
<position>299,-171</position>
<input>
<ID>IN_0</ID>64 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>296,-180.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>73 </input>
<input>
<ID>IN_2</ID>72 </input>
<input>
<ID>IN_3</ID>70 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_REGISTER4</type>
<position>287.5,-163.5</position>
<output>
<ID>OUT_0</ID>71 </output>
<output>
<ID>OUT_1</ID>73 </output>
<output>
<ID>OUT_2</ID>72 </output>
<output>
<ID>OUT_3</ID>70 </output>
<input>
<ID>clear</ID>74 </input>
<input>
<ID>clock</ID>68 </input>
<input>
<ID>count_enable</ID>68 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_AND2</type>
<position>288.5,-171</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>71 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>285.5,-180.5</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>78 </input>
<input>
<ID>IN_2</ID>77 </input>
<input>
<ID>IN_3</ID>75 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_REGISTER4</type>
<position>277,-163.5</position>
<output>
<ID>OUT_0</ID>76 </output>
<output>
<ID>OUT_1</ID>78 </output>
<output>
<ID>OUT_2</ID>77 </output>
<output>
<ID>OUT_3</ID>75 </output>
<input>
<ID>clear</ID>83 </input>
<input>
<ID>clock</ID>74 </input>
<input>
<ID>count_enable</ID>74 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>278,-171</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>275,-180.5</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>82 </input>
<input>
<ID>IN_2</ID>81 </input>
<input>
<ID>IN_3</ID>79 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_REGISTER4</type>
<position>266.5,-163.5</position>
<output>
<ID>OUT_0</ID>80 </output>
<output>
<ID>OUT_1</ID>82 </output>
<output>
<ID>OUT_2</ID>81 </output>
<output>
<ID>OUT_3</ID>79 </output>
<input>
<ID>clear</ID>89 </input>
<input>
<ID>clock</ID>83 </input>
<input>
<ID>count_enable</ID>83 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_AND2</type>
<position>267.5,-171</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>264.5,-180.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>87 </input>
<input>
<ID>IN_2</ID>86 </input>
<input>
<ID>IN_3</ID>84 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_REGISTER4</type>
<position>256,-163.5</position>
<output>
<ID>OUT_0</ID>85 </output>
<output>
<ID>OUT_1</ID>87 </output>
<output>
<ID>OUT_2</ID>86 </output>
<output>
<ID>OUT_3</ID>84 </output>
<input>
<ID>clear</ID>117 </input>
<input>
<ID>clock</ID>89 </input>
<input>
<ID>count_enable</ID>89 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_AND2</type>
<position>257,-171</position>
<input>
<ID>IN_0</ID>84 </input>
<input>
<ID>IN_1</ID>85 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>254,-180.5</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>94 </input>
<input>
<ID>IN_2</ID>93 </input>
<input>
<ID>IN_3</ID>91 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_REGISTER4</type>
<position>245.5,-163.5</position>
<output>
<ID>OUT_0</ID>92 </output>
<output>
<ID>OUT_1</ID>94 </output>
<output>
<ID>OUT_2</ID>93 </output>
<output>
<ID>OUT_3</ID>91 </output>
<input>
<ID>clear</ID>118 </input>
<input>
<ID>clock</ID>117 </input>
<input>
<ID>count_enable</ID>117 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_AND2</type>
<position>246.5,-171</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>92 </input>
<output>
<ID>OUT</ID>118 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>243.5,-180.5</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>99 </input>
<input>
<ID>IN_2</ID>98 </input>
<input>
<ID>IN_3</ID>96 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_REGISTER4</type>
<position>235,-163.5</position>
<output>
<ID>OUT_0</ID>97 </output>
<output>
<ID>OUT_1</ID>99 </output>
<output>
<ID>OUT_2</ID>98 </output>
<output>
<ID>OUT_3</ID>96 </output>
<input>
<ID>clear</ID>100 </input>
<input>
<ID>clock</ID>118 </input>
<input>
<ID>count_enable</ID>118 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_AND2</type>
<position>236,-171</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>233,-180.5</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>104 </input>
<input>
<ID>IN_2</ID>103 </input>
<input>
<ID>IN_3</ID>101 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_REGISTER4</type>
<position>224.5,-163.5</position>
<output>
<ID>OUT_0</ID>102 </output>
<output>
<ID>OUT_1</ID>104 </output>
<output>
<ID>OUT_2</ID>103 </output>
<output>
<ID>OUT_3</ID>101 </output>
<input>
<ID>clear</ID>109 </input>
<input>
<ID>clock</ID>100 </input>
<input>
<ID>count_enable</ID>100 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>59</ID>
<type>AA_AND2</type>
<position>225.5,-171</position>
<input>
<ID>IN_0</ID>101 </input>
<input>
<ID>IN_1</ID>102 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>222.5,-180.5</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>108 </input>
<input>
<ID>IN_2</ID>107 </input>
<input>
<ID>IN_3</ID>105 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_REGISTER4</type>
<position>214,-163.5</position>
<output>
<ID>OUT_0</ID>106 </output>
<output>
<ID>OUT_1</ID>108 </output>
<output>
<ID>OUT_2</ID>107 </output>
<output>
<ID>OUT_3</ID>105 </output>
<input>
<ID>clear</ID>115 </input>
<input>
<ID>clock</ID>109 </input>
<input>
<ID>count_enable</ID>109 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_AND2</type>
<position>215,-171</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>115 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>63</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>212,-180.5</position>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>113 </input>
<input>
<ID>IN_2</ID>112 </input>
<input>
<ID>IN_3</ID>110 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_REGISTER4</type>
<position>203.5,-163.5</position>
<output>
<ID>OUT_0</ID>111 </output>
<output>
<ID>OUT_1</ID>113 </output>
<output>
<ID>OUT_2</ID>112 </output>
<output>
<ID>OUT_3</ID>110 </output>
<input>
<ID>clear</ID>164 </input>
<input>
<ID>clock</ID>115 </input>
<input>
<ID>count_enable</ID>115 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_AND2</type>
<position>204.5,-171</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>111 </input>
<output>
<ID>OUT</ID>164 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_REGISTER4</type>
<position>266.5,-190</position>
<output>
<ID>OUT_0</ID>53 </output>
<output>
<ID>OUT_1</ID>55 </output>
<output>
<ID>OUT_2</ID>54 </output>
<output>
<ID>OUT_3</ID>52 </output>
<input>
<ID>clear</ID>61 </input>
<input>
<ID>clock</ID>56 </input>
<input>
<ID>count_enable</ID>56 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_AND2</type>
<position>267.5,-197.5</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>264.5,-207</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>60 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>57 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_REGISTER4</type>
<position>256,-190</position>
<output>
<ID>OUT_0</ID>58 </output>
<output>
<ID>OUT_1</ID>60 </output>
<output>
<ID>OUT_2</ID>59 </output>
<output>
<ID>OUT_3</ID>57 </output>
<input>
<ID>clear</ID>138 </input>
<input>
<ID>clock</ID>61 </input>
<input>
<ID>count_enable</ID>61 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_AND2</type>
<position>257,-197.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>58 </input>
<output>
<ID>OUT</ID>138 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>254,-207</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>95 </input>
<input>
<ID>IN_2</ID>88 </input>
<input>
<ID>IN_3</ID>63 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_REGISTER4</type>
<position>245.5,-190</position>
<output>
<ID>OUT_0</ID>69 </output>
<output>
<ID>OUT_1</ID>95 </output>
<output>
<ID>OUT_2</ID>88 </output>
<output>
<ID>OUT_3</ID>63 </output>
<input>
<ID>clear</ID>139 </input>
<input>
<ID>clock</ID>138 </input>
<input>
<ID>count_enable</ID>138 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_AND2</type>
<position>246.5,-197.5</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>139 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>243.5,-207</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>121 </input>
<input>
<ID>IN_2</ID>120 </input>
<input>
<ID>IN_3</ID>116 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_REGISTER4</type>
<position>235,-190</position>
<output>
<ID>OUT_0</ID>119 </output>
<output>
<ID>OUT_1</ID>121 </output>
<output>
<ID>OUT_2</ID>120 </output>
<output>
<ID>OUT_3</ID>116 </output>
<input>
<ID>clear</ID>122 </input>
<input>
<ID>clock</ID>139 </input>
<input>
<ID>count_enable</ID>139 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_AND2</type>
<position>236,-197.5</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>233,-207</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>126 </input>
<input>
<ID>IN_2</ID>125 </input>
<input>
<ID>IN_3</ID>123 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_REGISTER4</type>
<position>224.5,-190</position>
<output>
<ID>OUT_0</ID>124 </output>
<output>
<ID>OUT_1</ID>126 </output>
<output>
<ID>OUT_2</ID>125 </output>
<output>
<ID>OUT_3</ID>123 </output>
<input>
<ID>clear</ID>131 </input>
<input>
<ID>clock</ID>122 </input>
<input>
<ID>count_enable</ID>122 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_AND2</type>
<position>225.5,-197.5</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>131 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>222.5,-207</position>
<input>
<ID>IN_0</ID>128 </input>
<input>
<ID>IN_1</ID>130 </input>
<input>
<ID>IN_2</ID>129 </input>
<input>
<ID>IN_3</ID>127 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_REGISTER4</type>
<position>214,-190</position>
<output>
<ID>OUT_0</ID>128 </output>
<output>
<ID>OUT_1</ID>130 </output>
<output>
<ID>OUT_2</ID>129 </output>
<output>
<ID>OUT_3</ID>127 </output>
<input>
<ID>clear</ID>137 </input>
<input>
<ID>clock</ID>131 </input>
<input>
<ID>count_enable</ID>131 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_AND2</type>
<position>215,-197.5</position>
<input>
<ID>IN_0</ID>127 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>212,-207</position>
<input>
<ID>IN_0</ID>133 </input>
<input>
<ID>IN_1</ID>135 </input>
<input>
<ID>IN_2</ID>134 </input>
<input>
<ID>IN_3</ID>132 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_REGISTER4</type>
<position>203.5,-190</position>
<output>
<ID>OUT_0</ID>133 </output>
<output>
<ID>OUT_1</ID>135 </output>
<output>
<ID>OUT_2</ID>134 </output>
<output>
<ID>OUT_3</ID>132 </output>
<input>
<ID>clear</ID>90 </input>
<input>
<ID>clock</ID>137 </input>
<input>
<ID>count_enable</ID>137 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_AND2</type>
<position>204.5,-197.5</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>86</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>306,-153</position>
<input>
<ID>IN_0</ID>141 </input>
<input>
<ID>IN_1</ID>143 </input>
<input>
<ID>IN_2</ID>142 </input>
<input>
<ID>IN_3</ID>140 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>87</ID>
<type>AA_REGISTER4</type>
<position>297.5,-136</position>
<output>
<ID>OUT_0</ID>141 </output>
<output>
<ID>OUT_1</ID>143 </output>
<output>
<ID>OUT_2</ID>142 </output>
<output>
<ID>OUT_3</ID>140 </output>
<input>
<ID>clear</ID>144 </input>
<input>
<ID>clock</ID>164 </input>
<input>
<ID>count_enable</ID>164 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>88</ID>
<type>AA_AND2</type>
<position>298.5,-143.5</position>
<input>
<ID>IN_0</ID>140 </input>
<input>
<ID>IN_1</ID>141 </input>
<output>
<ID>OUT</ID>144 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>295.5,-153</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>148 </input>
<input>
<ID>IN_2</ID>147 </input>
<input>
<ID>IN_3</ID>145 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_REGISTER4</type>
<position>287,-136</position>
<output>
<ID>OUT_0</ID>146 </output>
<output>
<ID>OUT_1</ID>148 </output>
<output>
<ID>OUT_2</ID>147 </output>
<output>
<ID>OUT_3</ID>145 </output>
<input>
<ID>clear</ID>149 </input>
<input>
<ID>clock</ID>144 </input>
<input>
<ID>count_enable</ID>144 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>91</ID>
<type>AA_AND2</type>
<position>288,-143.5</position>
<input>
<ID>IN_0</ID>145 </input>
<input>
<ID>IN_1</ID>146 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>285,-153</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>153 </input>
<input>
<ID>IN_2</ID>152 </input>
<input>
<ID>IN_3</ID>150 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>93</ID>
<type>AA_REGISTER4</type>
<position>276.5,-136</position>
<output>
<ID>OUT_0</ID>151 </output>
<output>
<ID>OUT_1</ID>153 </output>
<output>
<ID>OUT_2</ID>152 </output>
<output>
<ID>OUT_3</ID>150 </output>
<input>
<ID>clear</ID>158 </input>
<input>
<ID>clock</ID>149 </input>
<input>
<ID>count_enable</ID>149 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_AND2</type>
<position>277.5,-143.5</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>151 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>274.5,-153</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>157 </input>
<input>
<ID>IN_2</ID>156 </input>
<input>
<ID>IN_3</ID>154 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>96</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>306,-126.5</position>
<input>
<ID>IN_0</ID>167 </input>
<input>
<ID>IN_1</ID>169 </input>
<input>
<ID>IN_2</ID>168 </input>
<input>
<ID>IN_3</ID>166 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_REGISTER4</type>
<position>297.5,-109.5</position>
<output>
<ID>OUT_0</ID>167 </output>
<output>
<ID>OUT_1</ID>169 </output>
<output>
<ID>OUT_2</ID>168 </output>
<output>
<ID>OUT_3</ID>166 </output>
<input>
<ID>clear</ID>170 </input>
<input>
<ID>clock</ID>192 </input>
<input>
<ID>count_enable</ID>192 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_AND2</type>
<position>298.5,-117</position>
<input>
<ID>IN_0</ID>166 </input>
<input>
<ID>IN_1</ID>167 </input>
<output>
<ID>OUT</ID>170 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>295.5,-126.5</position>
<input>
<ID>IN_0</ID>173 </input>
<input>
<ID>IN_1</ID>175 </input>
<input>
<ID>IN_2</ID>174 </input>
<input>
<ID>IN_3</ID>172 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>100</ID>
<type>AA_REGISTER4</type>
<position>287,-109.5</position>
<output>
<ID>OUT_0</ID>173 </output>
<output>
<ID>OUT_1</ID>175 </output>
<output>
<ID>OUT_2</ID>174 </output>
<output>
<ID>OUT_3</ID>172 </output>
<input>
<ID>clear</ID>176 </input>
<input>
<ID>clock</ID>170 </input>
<input>
<ID>count_enable</ID>170 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_AND2</type>
<position>288,-117</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>173 </input>
<output>
<ID>OUT</ID>176 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>285,-126.5</position>
<input>
<ID>IN_0</ID>178 </input>
<input>
<ID>IN_1</ID>180 </input>
<input>
<ID>IN_2</ID>179 </input>
<input>
<ID>IN_3</ID>177 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_REGISTER4</type>
<position>276.5,-109.5</position>
<output>
<ID>OUT_0</ID>178 </output>
<output>
<ID>OUT_1</ID>180 </output>
<output>
<ID>OUT_2</ID>179 </output>
<output>
<ID>OUT_3</ID>177 </output>
<input>
<ID>clear</ID>185 </input>
<input>
<ID>clock</ID>176 </input>
<input>
<ID>count_enable</ID>176 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_AND2</type>
<position>277.5,-117</position>
<input>
<ID>IN_0</ID>177 </input>
<input>
<ID>IN_1</ID>178 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>105</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>274.5,-126.5</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>184 </input>
<input>
<ID>IN_2</ID>183 </input>
<input>
<ID>IN_3</ID>181 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_REGISTER4</type>
<position>266,-109.5</position>
<output>
<ID>OUT_0</ID>182 </output>
<output>
<ID>OUT_1</ID>184 </output>
<output>
<ID>OUT_2</ID>183 </output>
<output>
<ID>OUT_3</ID>181 </output>
<input>
<ID>clear</ID>191 </input>
<input>
<ID>clock</ID>185 </input>
<input>
<ID>count_enable</ID>185 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_AND2</type>
<position>267,-117</position>
<input>
<ID>IN_0</ID>181 </input>
<input>
<ID>IN_1</ID>182 </input>
<output>
<ID>OUT</ID>191 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>264,-126.5</position>
<input>
<ID>IN_0</ID>187 </input>
<input>
<ID>IN_1</ID>189 </input>
<input>
<ID>IN_2</ID>188 </input>
<input>
<ID>IN_3</ID>186 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_REGISTER4</type>
<position>255.5,-109.5</position>
<output>
<ID>OUT_0</ID>187 </output>
<output>
<ID>OUT_1</ID>189 </output>
<output>
<ID>OUT_2</ID>188 </output>
<output>
<ID>OUT_3</ID>186 </output>
<input>
<ID>clear</ID>219 </input>
<input>
<ID>clock</ID>191 </input>
<input>
<ID>count_enable</ID>191 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_AND2</type>
<position>256.5,-117</position>
<input>
<ID>IN_0</ID>186 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>219 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>111</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>253.5,-126.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>196 </input>
<input>
<ID>IN_2</ID>195 </input>
<input>
<ID>IN_3</ID>193 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_REGISTER4</type>
<position>245,-109.5</position>
<output>
<ID>OUT_0</ID>194 </output>
<output>
<ID>OUT_1</ID>196 </output>
<output>
<ID>OUT_2</ID>195 </output>
<output>
<ID>OUT_3</ID>193 </output>
<input>
<ID>clear</ID>220 </input>
<input>
<ID>clock</ID>219 </input>
<input>
<ID>count_enable</ID>219 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_AND2</type>
<position>246,-117</position>
<input>
<ID>IN_0</ID>193 </input>
<input>
<ID>IN_1</ID>194 </input>
<output>
<ID>OUT</ID>220 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>243,-126.5</position>
<input>
<ID>IN_0</ID>199 </input>
<input>
<ID>IN_1</ID>201 </input>
<input>
<ID>IN_2</ID>200 </input>
<input>
<ID>IN_3</ID>198 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_REGISTER4</type>
<position>234.5,-109.5</position>
<output>
<ID>OUT_0</ID>199 </output>
<output>
<ID>OUT_1</ID>201 </output>
<output>
<ID>OUT_2</ID>200 </output>
<output>
<ID>OUT_3</ID>198 </output>
<input>
<ID>clear</ID>202 </input>
<input>
<ID>clock</ID>220 </input>
<input>
<ID>count_enable</ID>220 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_AND2</type>
<position>235.5,-117</position>
<input>
<ID>IN_0</ID>198 </input>
<input>
<ID>IN_1</ID>199 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>232.5,-126.5</position>
<input>
<ID>IN_0</ID>204 </input>
<input>
<ID>IN_1</ID>206 </input>
<input>
<ID>IN_2</ID>205 </input>
<input>
<ID>IN_3</ID>203 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>118</ID>
<type>AA_REGISTER4</type>
<position>224,-109.5</position>
<output>
<ID>OUT_0</ID>204 </output>
<output>
<ID>OUT_1</ID>206 </output>
<output>
<ID>OUT_2</ID>205 </output>
<output>
<ID>OUT_3</ID>203 </output>
<input>
<ID>clear</ID>211 </input>
<input>
<ID>clock</ID>202 </input>
<input>
<ID>count_enable</ID>202 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_AND2</type>
<position>225,-117</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>204 </input>
<output>
<ID>OUT</ID>211 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>222,-126.5</position>
<input>
<ID>IN_0</ID>208 </input>
<input>
<ID>IN_1</ID>210 </input>
<input>
<ID>IN_2</ID>209 </input>
<input>
<ID>IN_3</ID>207 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_REGISTER4</type>
<position>213.5,-109.5</position>
<output>
<ID>OUT_0</ID>208 </output>
<output>
<ID>OUT_1</ID>210 </output>
<output>
<ID>OUT_2</ID>209 </output>
<output>
<ID>OUT_3</ID>207 </output>
<input>
<ID>clear</ID>217 </input>
<input>
<ID>clock</ID>211 </input>
<input>
<ID>count_enable</ID>211 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_AND2</type>
<position>214.5,-117</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>211.5,-126.5</position>
<input>
<ID>IN_0</ID>213 </input>
<input>
<ID>IN_1</ID>215 </input>
<input>
<ID>IN_2</ID>214 </input>
<input>
<ID>IN_3</ID>212 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_REGISTER4</type>
<position>203,-109.5</position>
<output>
<ID>OUT_0</ID>213 </output>
<output>
<ID>OUT_1</ID>215 </output>
<output>
<ID>OUT_2</ID>214 </output>
<output>
<ID>OUT_3</ID>212 </output>
<input>
<ID>clear</ID>265 </input>
<input>
<ID>clock</ID>217 </input>
<input>
<ID>count_enable</ID>217 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_AND2</type>
<position>204,-117</position>
<input>
<ID>IN_0</ID>212 </input>
<input>
<ID>IN_1</ID>213 </input>
<output>
<ID>OUT</ID>265 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_REGISTER4</type>
<position>266,-136</position>
<output>
<ID>OUT_0</ID>155 </output>
<output>
<ID>OUT_1</ID>157 </output>
<output>
<ID>OUT_2</ID>156 </output>
<output>
<ID>OUT_3</ID>154 </output>
<input>
<ID>clear</ID>163 </input>
<input>
<ID>clock</ID>158 </input>
<input>
<ID>count_enable</ID>158 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_AND2</type>
<position>267,-143.5</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>155 </input>
<output>
<ID>OUT</ID>163 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>128</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>264,-153</position>
<input>
<ID>IN_0</ID>160 </input>
<input>
<ID>IN_1</ID>162 </input>
<input>
<ID>IN_2</ID>161 </input>
<input>
<ID>IN_3</ID>159 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>129</ID>
<type>AA_REGISTER4</type>
<position>255.5,-136</position>
<output>
<ID>OUT_0</ID>160 </output>
<output>
<ID>OUT_1</ID>162 </output>
<output>
<ID>OUT_2</ID>161 </output>
<output>
<ID>OUT_3</ID>159 </output>
<input>
<ID>clear</ID>239 </input>
<input>
<ID>clock</ID>163 </input>
<input>
<ID>count_enable</ID>163 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_AND2</type>
<position>256.5,-143.5</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>160 </input>
<output>
<ID>OUT</ID>239 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>131</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>253.5,-153</position>
<input>
<ID>IN_0</ID>171 </input>
<input>
<ID>IN_1</ID>197 </input>
<input>
<ID>IN_2</ID>190 </input>
<input>
<ID>IN_3</ID>165 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_REGISTER4</type>
<position>245,-136</position>
<output>
<ID>OUT_0</ID>171 </output>
<output>
<ID>OUT_1</ID>197 </output>
<output>
<ID>OUT_2</ID>190 </output>
<output>
<ID>OUT_3</ID>165 </output>
<input>
<ID>clear</ID>240 </input>
<input>
<ID>clock</ID>239 </input>
<input>
<ID>count_enable</ID>239 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>133</ID>
<type>AA_AND2</type>
<position>246,-143.5</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>171 </input>
<output>
<ID>OUT</ID>240 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>243,-153</position>
<input>
<ID>IN_0</ID>221 </input>
<input>
<ID>IN_1</ID>223 </input>
<input>
<ID>IN_2</ID>222 </input>
<input>
<ID>IN_3</ID>218 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>135</ID>
<type>AA_REGISTER4</type>
<position>234.5,-136</position>
<output>
<ID>OUT_0</ID>221 </output>
<output>
<ID>OUT_1</ID>223 </output>
<output>
<ID>OUT_2</ID>222 </output>
<output>
<ID>OUT_3</ID>218 </output>
<input>
<ID>clear</ID>224 </input>
<input>
<ID>clock</ID>240 </input>
<input>
<ID>count_enable</ID>240 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>136</ID>
<type>AA_AND2</type>
<position>235.5,-143.5</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>221 </input>
<output>
<ID>OUT</ID>224 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>137</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>232.5,-153</position>
<input>
<ID>IN_0</ID>226 </input>
<input>
<ID>IN_1</ID>228 </input>
<input>
<ID>IN_2</ID>227 </input>
<input>
<ID>IN_3</ID>225 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_REGISTER4</type>
<position>224,-136</position>
<output>
<ID>OUT_0</ID>226 </output>
<output>
<ID>OUT_1</ID>228 </output>
<output>
<ID>OUT_2</ID>227 </output>
<output>
<ID>OUT_3</ID>225 </output>
<input>
<ID>clear</ID>233 </input>
<input>
<ID>clock</ID>224 </input>
<input>
<ID>count_enable</ID>224 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>139</ID>
<type>AA_AND2</type>
<position>225,-143.5</position>
<input>
<ID>IN_0</ID>225 </input>
<input>
<ID>IN_1</ID>226 </input>
<output>
<ID>OUT</ID>233 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>140</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>222,-153</position>
<input>
<ID>IN_0</ID>230 </input>
<input>
<ID>IN_1</ID>232 </input>
<input>
<ID>IN_2</ID>231 </input>
<input>
<ID>IN_3</ID>229 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_REGISTER4</type>
<position>213.5,-136</position>
<output>
<ID>OUT_0</ID>230 </output>
<output>
<ID>OUT_1</ID>232 </output>
<output>
<ID>OUT_2</ID>231 </output>
<output>
<ID>OUT_3</ID>229 </output>
<input>
<ID>clear</ID>238 </input>
<input>
<ID>clock</ID>233 </input>
<input>
<ID>count_enable</ID>233 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_AND2</type>
<position>214.5,-143.5</position>
<input>
<ID>IN_0</ID>229 </input>
<input>
<ID>IN_1</ID>230 </input>
<output>
<ID>OUT</ID>238 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>143</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>211.5,-153</position>
<input>
<ID>IN_0</ID>235 </input>
<input>
<ID>IN_1</ID>237 </input>
<input>
<ID>IN_2</ID>236 </input>
<input>
<ID>IN_3</ID>234 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_REGISTER4</type>
<position>203,-136</position>
<output>
<ID>OUT_0</ID>235 </output>
<output>
<ID>OUT_1</ID>237 </output>
<output>
<ID>OUT_2</ID>236 </output>
<output>
<ID>OUT_3</ID>234 </output>
<input>
<ID>clear</ID>192 </input>
<input>
<ID>clock</ID>238 </input>
<input>
<ID>count_enable</ID>238 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_AND2</type>
<position>204,-143.5</position>
<input>
<ID>IN_0</ID>234 </input>
<input>
<ID>IN_1</ID>235 </input>
<output>
<ID>OUT</ID>192 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>146</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>306,-99</position>
<input>
<ID>IN_0</ID>242 </input>
<input>
<ID>IN_1</ID>244 </input>
<input>
<ID>IN_2</ID>243 </input>
<input>
<ID>IN_3</ID>241 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_REGISTER4</type>
<position>297.5,-82</position>
<output>
<ID>OUT_0</ID>242 </output>
<output>
<ID>OUT_1</ID>244 </output>
<output>
<ID>OUT_2</ID>243 </output>
<output>
<ID>OUT_3</ID>241 </output>
<input>
<ID>clear</ID>245 </input>
<input>
<ID>clock</ID>265 </input>
<input>
<ID>count_enable</ID>265 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>148</ID>
<type>AA_AND2</type>
<position>298.5,-89.5</position>
<input>
<ID>IN_0</ID>241 </input>
<input>
<ID>IN_1</ID>242 </input>
<output>
<ID>OUT</ID>245 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>149</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>295.5,-99</position>
<input>
<ID>IN_0</ID>247 </input>
<input>
<ID>IN_1</ID>249 </input>
<input>
<ID>IN_2</ID>248 </input>
<input>
<ID>IN_3</ID>246 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_REGISTER4</type>
<position>287,-82</position>
<output>
<ID>OUT_0</ID>247 </output>
<output>
<ID>OUT_1</ID>249 </output>
<output>
<ID>OUT_2</ID>248 </output>
<output>
<ID>OUT_3</ID>246 </output>
<input>
<ID>clear</ID>250 </input>
<input>
<ID>clock</ID>245 </input>
<input>
<ID>count_enable</ID>245 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_AND2</type>
<position>288,-89.5</position>
<input>
<ID>IN_0</ID>246 </input>
<input>
<ID>IN_1</ID>247 </input>
<output>
<ID>OUT</ID>250 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>152</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>285,-99</position>
<input>
<ID>IN_0</ID>252 </input>
<input>
<ID>IN_1</ID>254 </input>
<input>
<ID>IN_2</ID>253 </input>
<input>
<ID>IN_3</ID>251 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_REGISTER4</type>
<position>276.5,-82</position>
<output>
<ID>OUT_0</ID>252 </output>
<output>
<ID>OUT_1</ID>254 </output>
<output>
<ID>OUT_2</ID>253 </output>
<output>
<ID>OUT_3</ID>251 </output>
<input>
<ID>clear</ID>259 </input>
<input>
<ID>clock</ID>250 </input>
<input>
<ID>count_enable</ID>250 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>154</ID>
<type>AA_AND2</type>
<position>277.5,-89.5</position>
<input>
<ID>IN_0</ID>251 </input>
<input>
<ID>IN_1</ID>252 </input>
<output>
<ID>OUT</ID>259 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>155</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>274.5,-99</position>
<input>
<ID>IN_0</ID>256 </input>
<input>
<ID>IN_1</ID>258 </input>
<input>
<ID>IN_2</ID>257 </input>
<input>
<ID>IN_3</ID>255 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>156</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>306,-72.5</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>270 </input>
<input>
<ID>IN_2</ID>269 </input>
<input>
<ID>IN_3</ID>267 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_REGISTER4</type>
<position>297.5,-55.5</position>
<output>
<ID>OUT_0</ID>268 </output>
<output>
<ID>OUT_1</ID>270 </output>
<output>
<ID>OUT_2</ID>269 </output>
<output>
<ID>OUT_3</ID>267 </output>
<input>
<ID>clear</ID>271 </input>
<input>
<ID>clock</ID>293 </input>
<input>
<ID>count_enable</ID>293 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>158</ID>
<type>AA_AND2</type>
<position>298.5,-63</position>
<input>
<ID>IN_0</ID>267 </input>
<input>
<ID>IN_1</ID>268 </input>
<output>
<ID>OUT</ID>271 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>159</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>295.5,-72.5</position>
<input>
<ID>IN_0</ID>274 </input>
<input>
<ID>IN_1</ID>276 </input>
<input>
<ID>IN_2</ID>275 </input>
<input>
<ID>IN_3</ID>273 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>160</ID>
<type>AA_REGISTER4</type>
<position>287,-55.5</position>
<output>
<ID>OUT_0</ID>274 </output>
<output>
<ID>OUT_1</ID>276 </output>
<output>
<ID>OUT_2</ID>275 </output>
<output>
<ID>OUT_3</ID>273 </output>
<input>
<ID>clear</ID>277 </input>
<input>
<ID>clock</ID>271 </input>
<input>
<ID>count_enable</ID>271 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_AND2</type>
<position>288,-63</position>
<input>
<ID>IN_0</ID>273 </input>
<input>
<ID>IN_1</ID>274 </input>
<output>
<ID>OUT</ID>277 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>162</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>285,-72.5</position>
<input>
<ID>IN_0</ID>279 </input>
<input>
<ID>IN_1</ID>281 </input>
<input>
<ID>IN_2</ID>280 </input>
<input>
<ID>IN_3</ID>278 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>163</ID>
<type>AA_REGISTER4</type>
<position>276.5,-55.5</position>
<output>
<ID>OUT_0</ID>279 </output>
<output>
<ID>OUT_1</ID>281 </output>
<output>
<ID>OUT_2</ID>280 </output>
<output>
<ID>OUT_3</ID>278 </output>
<input>
<ID>clear</ID>286 </input>
<input>
<ID>clock</ID>277 </input>
<input>
<ID>count_enable</ID>277 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>164</ID>
<type>AA_AND2</type>
<position>277.5,-63</position>
<input>
<ID>IN_0</ID>278 </input>
<input>
<ID>IN_1</ID>279 </input>
<output>
<ID>OUT</ID>286 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>165</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>274.5,-72.5</position>
<input>
<ID>IN_0</ID>283 </input>
<input>
<ID>IN_1</ID>285 </input>
<input>
<ID>IN_2</ID>284 </input>
<input>
<ID>IN_3</ID>282 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>166</ID>
<type>AA_REGISTER4</type>
<position>266,-55.5</position>
<output>
<ID>OUT_0</ID>283 </output>
<output>
<ID>OUT_1</ID>285 </output>
<output>
<ID>OUT_2</ID>284 </output>
<output>
<ID>OUT_3</ID>282 </output>
<input>
<ID>clear</ID>292 </input>
<input>
<ID>clock</ID>286 </input>
<input>
<ID>count_enable</ID>286 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_AND2</type>
<position>267,-63</position>
<input>
<ID>IN_0</ID>282 </input>
<input>
<ID>IN_1</ID>283 </input>
<output>
<ID>OUT</ID>292 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>168</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>264,-72.5</position>
<input>
<ID>IN_0</ID>288 </input>
<input>
<ID>IN_1</ID>290 </input>
<input>
<ID>IN_2</ID>289 </input>
<input>
<ID>IN_3</ID>287 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_REGISTER4</type>
<position>255.5,-55.5</position>
<output>
<ID>OUT_0</ID>288 </output>
<output>
<ID>OUT_1</ID>290 </output>
<output>
<ID>OUT_2</ID>289 </output>
<output>
<ID>OUT_3</ID>287 </output>
<input>
<ID>clear</ID>319 </input>
<input>
<ID>clock</ID>292 </input>
<input>
<ID>count_enable</ID>292 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_AND2</type>
<position>256.5,-63</position>
<input>
<ID>IN_0</ID>287 </input>
<input>
<ID>IN_1</ID>288 </input>
<output>
<ID>OUT</ID>319 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>171</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>253.5,-72.5</position>
<input>
<ID>IN_0</ID>295 </input>
<input>
<ID>IN_1</ID>297 </input>
<input>
<ID>IN_2</ID>296 </input>
<input>
<ID>IN_3</ID>294 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_REGISTER4</type>
<position>245,-55.5</position>
<output>
<ID>OUT_0</ID>295 </output>
<output>
<ID>OUT_1</ID>297 </output>
<output>
<ID>OUT_2</ID>296 </output>
<output>
<ID>OUT_3</ID>294 </output>
<input>
<ID>clear</ID>320 </input>
<input>
<ID>clock</ID>319 </input>
<input>
<ID>count_enable</ID>319 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_AND2</type>
<position>246,-63</position>
<input>
<ID>IN_0</ID>294 </input>
<input>
<ID>IN_1</ID>295 </input>
<output>
<ID>OUT</ID>320 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>174</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>243,-72.5</position>
<input>
<ID>IN_0</ID>300 </input>
<input>
<ID>IN_1</ID>302 </input>
<input>
<ID>IN_2</ID>301 </input>
<input>
<ID>IN_3</ID>299 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>175</ID>
<type>AA_REGISTER4</type>
<position>234.5,-55.5</position>
<output>
<ID>OUT_0</ID>300 </output>
<output>
<ID>OUT_1</ID>302 </output>
<output>
<ID>OUT_2</ID>301 </output>
<output>
<ID>OUT_3</ID>299 </output>
<input>
<ID>clear</ID>303 </input>
<input>
<ID>clock</ID>320 </input>
<input>
<ID>count_enable</ID>320 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_AND2</type>
<position>235.5,-63</position>
<input>
<ID>IN_0</ID>299 </input>
<input>
<ID>IN_1</ID>300 </input>
<output>
<ID>OUT</ID>303 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>232.5,-72.5</position>
<input>
<ID>IN_0</ID>305 </input>
<input>
<ID>IN_1</ID>307 </input>
<input>
<ID>IN_2</ID>306 </input>
<input>
<ID>IN_3</ID>304 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_REGISTER4</type>
<position>224,-55.5</position>
<output>
<ID>OUT_0</ID>305 </output>
<output>
<ID>OUT_1</ID>307 </output>
<output>
<ID>OUT_2</ID>306 </output>
<output>
<ID>OUT_3</ID>304 </output>
<input>
<ID>clear</ID>312 </input>
<input>
<ID>clock</ID>303 </input>
<input>
<ID>count_enable</ID>303 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_AND2</type>
<position>225,-63</position>
<input>
<ID>IN_0</ID>304 </input>
<input>
<ID>IN_1</ID>305 </input>
<output>
<ID>OUT</ID>312 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>180</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>222,-72.5</position>
<input>
<ID>IN_0</ID>309 </input>
<input>
<ID>IN_1</ID>311 </input>
<input>
<ID>IN_2</ID>310 </input>
<input>
<ID>IN_3</ID>308 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_REGISTER4</type>
<position>213.5,-55.5</position>
<output>
<ID>OUT_0</ID>309 </output>
<output>
<ID>OUT_1</ID>311 </output>
<output>
<ID>OUT_2</ID>310 </output>
<output>
<ID>OUT_3</ID>308 </output>
<input>
<ID>clear</ID>317 </input>
<input>
<ID>clock</ID>312 </input>
<input>
<ID>count_enable</ID>312 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_AND2</type>
<position>214.5,-63</position>
<input>
<ID>IN_0</ID>308 </input>
<input>
<ID>IN_1</ID>309 </input>
<output>
<ID>OUT</ID>317 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>183</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>211.5,-72.5</position>
<input>
<ID>IN_0</ID>314 </input>
<input>
<ID>IN_1</ID>316 </input>
<input>
<ID>IN_2</ID>315 </input>
<input>
<ID>IN_3</ID>313 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_REGISTER4</type>
<position>203,-55.5</position>
<output>
<ID>OUT_0</ID>314 </output>
<output>
<ID>OUT_1</ID>316 </output>
<output>
<ID>OUT_2</ID>315 </output>
<output>
<ID>OUT_3</ID>313 </output>
<input>
<ID>clear</ID>365 </input>
<input>
<ID>clock</ID>317 </input>
<input>
<ID>count_enable</ID>317 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>185</ID>
<type>AA_AND2</type>
<position>204,-63</position>
<input>
<ID>IN_0</ID>313 </input>
<input>
<ID>IN_1</ID>314 </input>
<output>
<ID>OUT</ID>365 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>186</ID>
<type>AA_REGISTER4</type>
<position>266,-82</position>
<output>
<ID>OUT_0</ID>256 </output>
<output>
<ID>OUT_1</ID>258 </output>
<output>
<ID>OUT_2</ID>257 </output>
<output>
<ID>OUT_3</ID>255 </output>
<input>
<ID>clear</ID>264 </input>
<input>
<ID>clock</ID>259 </input>
<input>
<ID>count_enable</ID>259 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>187</ID>
<type>AA_AND2</type>
<position>267,-89.5</position>
<input>
<ID>IN_0</ID>255 </input>
<input>
<ID>IN_1</ID>256 </input>
<output>
<ID>OUT</ID>264 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>188</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>264,-99</position>
<input>
<ID>IN_0</ID>261 </input>
<input>
<ID>IN_1</ID>263 </input>
<input>
<ID>IN_2</ID>262 </input>
<input>
<ID>IN_3</ID>260 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>189</ID>
<type>AA_REGISTER4</type>
<position>255.5,-82</position>
<output>
<ID>OUT_0</ID>261 </output>
<output>
<ID>OUT_1</ID>263 </output>
<output>
<ID>OUT_2</ID>262 </output>
<output>
<ID>OUT_3</ID>260 </output>
<input>
<ID>clear</ID>339 </input>
<input>
<ID>clock</ID>264 </input>
<input>
<ID>count_enable</ID>264 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_AND2</type>
<position>256.5,-89.5</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>261 </input>
<output>
<ID>OUT</ID>339 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>191</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>253.5,-99</position>
<input>
<ID>IN_0</ID>272 </input>
<input>
<ID>IN_1</ID>298 </input>
<input>
<ID>IN_2</ID>291 </input>
<input>
<ID>IN_3</ID>266 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_REGISTER4</type>
<position>245,-82</position>
<output>
<ID>OUT_0</ID>272 </output>
<output>
<ID>OUT_1</ID>298 </output>
<output>
<ID>OUT_2</ID>291 </output>
<output>
<ID>OUT_3</ID>266 </output>
<input>
<ID>clear</ID>340 </input>
<input>
<ID>clock</ID>339 </input>
<input>
<ID>count_enable</ID>339 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>193</ID>
<type>AA_AND2</type>
<position>246,-89.5</position>
<input>
<ID>IN_0</ID>266 </input>
<input>
<ID>IN_1</ID>272 </input>
<output>
<ID>OUT</ID>340 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>194</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>243,-99</position>
<input>
<ID>IN_0</ID>321 </input>
<input>
<ID>IN_1</ID>323 </input>
<input>
<ID>IN_2</ID>322 </input>
<input>
<ID>IN_3</ID>318 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>195</ID>
<type>AA_REGISTER4</type>
<position>234.5,-82</position>
<output>
<ID>OUT_0</ID>321 </output>
<output>
<ID>OUT_1</ID>323 </output>
<output>
<ID>OUT_2</ID>322 </output>
<output>
<ID>OUT_3</ID>318 </output>
<input>
<ID>clear</ID>324 </input>
<input>
<ID>clock</ID>340 </input>
<input>
<ID>count_enable</ID>340 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>196</ID>
<type>AA_AND2</type>
<position>235.5,-89.5</position>
<input>
<ID>IN_0</ID>318 </input>
<input>
<ID>IN_1</ID>321 </input>
<output>
<ID>OUT</ID>324 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>197</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>232.5,-99</position>
<input>
<ID>IN_0</ID>326 </input>
<input>
<ID>IN_1</ID>328 </input>
<input>
<ID>IN_2</ID>327 </input>
<input>
<ID>IN_3</ID>325 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_REGISTER4</type>
<position>224,-82</position>
<output>
<ID>OUT_0</ID>326 </output>
<output>
<ID>OUT_1</ID>328 </output>
<output>
<ID>OUT_2</ID>327 </output>
<output>
<ID>OUT_3</ID>325 </output>
<input>
<ID>clear</ID>333 </input>
<input>
<ID>clock</ID>324 </input>
<input>
<ID>count_enable</ID>324 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>199</ID>
<type>AA_AND2</type>
<position>225,-89.5</position>
<input>
<ID>IN_0</ID>325 </input>
<input>
<ID>IN_1</ID>326 </input>
<output>
<ID>OUT</ID>333 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>200</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>222,-99</position>
<input>
<ID>IN_0</ID>330 </input>
<input>
<ID>IN_1</ID>332 </input>
<input>
<ID>IN_2</ID>331 </input>
<input>
<ID>IN_3</ID>329 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_REGISTER4</type>
<position>213.5,-82</position>
<output>
<ID>OUT_0</ID>330 </output>
<output>
<ID>OUT_1</ID>332 </output>
<output>
<ID>OUT_2</ID>331 </output>
<output>
<ID>OUT_3</ID>329 </output>
<input>
<ID>clear</ID>338 </input>
<input>
<ID>clock</ID>333 </input>
<input>
<ID>count_enable</ID>333 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>202</ID>
<type>AA_AND2</type>
<position>214.5,-89.5</position>
<input>
<ID>IN_0</ID>329 </input>
<input>
<ID>IN_1</ID>330 </input>
<output>
<ID>OUT</ID>338 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>203</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>211.5,-99</position>
<input>
<ID>IN_0</ID>335 </input>
<input>
<ID>IN_1</ID>337 </input>
<input>
<ID>IN_2</ID>336 </input>
<input>
<ID>IN_3</ID>334 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>204</ID>
<type>AA_REGISTER4</type>
<position>203,-82</position>
<output>
<ID>OUT_0</ID>335 </output>
<output>
<ID>OUT_1</ID>337 </output>
<output>
<ID>OUT_2</ID>336 </output>
<output>
<ID>OUT_3</ID>334 </output>
<input>
<ID>clear</ID>293 </input>
<input>
<ID>clock</ID>338 </input>
<input>
<ID>count_enable</ID>338 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>205</ID>
<type>AA_AND2</type>
<position>204,-89.5</position>
<input>
<ID>IN_0</ID>334 </input>
<input>
<ID>IN_1</ID>335 </input>
<output>
<ID>OUT</ID>293 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>206</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>305.5,-45</position>
<input>
<ID>IN_0</ID>342 </input>
<input>
<ID>IN_1</ID>344 </input>
<input>
<ID>IN_2</ID>343 </input>
<input>
<ID>IN_3</ID>341 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>207</ID>
<type>AA_REGISTER4</type>
<position>297,-28</position>
<output>
<ID>OUT_0</ID>342 </output>
<output>
<ID>OUT_1</ID>344 </output>
<output>
<ID>OUT_2</ID>343 </output>
<output>
<ID>OUT_3</ID>341 </output>
<input>
<ID>clear</ID>345 </input>
<input>
<ID>clock</ID>365 </input>
<input>
<ID>count_enable</ID>365 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>208</ID>
<type>AA_AND2</type>
<position>298,-35.5</position>
<input>
<ID>IN_0</ID>341 </input>
<input>
<ID>IN_1</ID>342 </input>
<output>
<ID>OUT</ID>345 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>209</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>295,-45</position>
<input>
<ID>IN_0</ID>347 </input>
<input>
<ID>IN_1</ID>349 </input>
<input>
<ID>IN_2</ID>348 </input>
<input>
<ID>IN_3</ID>346 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>210</ID>
<type>AA_REGISTER4</type>
<position>286.5,-28</position>
<output>
<ID>OUT_0</ID>347 </output>
<output>
<ID>OUT_1</ID>349 </output>
<output>
<ID>OUT_2</ID>348 </output>
<output>
<ID>OUT_3</ID>346 </output>
<input>
<ID>clear</ID>350 </input>
<input>
<ID>clock</ID>345 </input>
<input>
<ID>count_enable</ID>345 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>211</ID>
<type>AA_AND2</type>
<position>287.5,-35.5</position>
<input>
<ID>IN_0</ID>346 </input>
<input>
<ID>IN_1</ID>347 </input>
<output>
<ID>OUT</ID>350 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>212</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>284.5,-45</position>
<input>
<ID>IN_0</ID>352 </input>
<input>
<ID>IN_1</ID>354 </input>
<input>
<ID>IN_2</ID>353 </input>
<input>
<ID>IN_3</ID>351 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>213</ID>
<type>AA_REGISTER4</type>
<position>276,-28</position>
<output>
<ID>OUT_0</ID>352 </output>
<output>
<ID>OUT_1</ID>354 </output>
<output>
<ID>OUT_2</ID>353 </output>
<output>
<ID>OUT_3</ID>351 </output>
<input>
<ID>clear</ID>359 </input>
<input>
<ID>clock</ID>350 </input>
<input>
<ID>count_enable</ID>350 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_AND2</type>
<position>277,-35.5</position>
<input>
<ID>IN_0</ID>351 </input>
<input>
<ID>IN_1</ID>352 </input>
<output>
<ID>OUT</ID>359 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>274,-45</position>
<input>
<ID>IN_0</ID>356 </input>
<input>
<ID>IN_1</ID>358 </input>
<input>
<ID>IN_2</ID>357 </input>
<input>
<ID>IN_3</ID>355 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>216</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>305.5,-18.5</position>
<input>
<ID>IN_0</ID>368 </input>
<input>
<ID>IN_1</ID>370 </input>
<input>
<ID>IN_2</ID>369 </input>
<input>
<ID>IN_3</ID>367 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>217</ID>
<type>AA_REGISTER4</type>
<position>297,-1.5</position>
<output>
<ID>OUT_0</ID>368 </output>
<output>
<ID>OUT_1</ID>370 </output>
<output>
<ID>OUT_2</ID>369 </output>
<output>
<ID>OUT_3</ID>367 </output>
<input>
<ID>clear</ID>371 </input>
<input>
<ID>clock</ID>393 </input>
<input>
<ID>count_enable</ID>393 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>218</ID>
<type>AA_AND2</type>
<position>298,-9</position>
<input>
<ID>IN_0</ID>367 </input>
<input>
<ID>IN_1</ID>368 </input>
<output>
<ID>OUT</ID>371 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>219</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>295,-18.5</position>
<input>
<ID>IN_0</ID>374 </input>
<input>
<ID>IN_1</ID>376 </input>
<input>
<ID>IN_2</ID>375 </input>
<input>
<ID>IN_3</ID>373 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_REGISTER4</type>
<position>286.5,-1.5</position>
<output>
<ID>OUT_0</ID>374 </output>
<output>
<ID>OUT_1</ID>376 </output>
<output>
<ID>OUT_2</ID>375 </output>
<output>
<ID>OUT_3</ID>373 </output>
<input>
<ID>clear</ID>377 </input>
<input>
<ID>clock</ID>371 </input>
<input>
<ID>count_enable</ID>371 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_AND2</type>
<position>287.5,-9</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>374 </input>
<output>
<ID>OUT</ID>377 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>284.5,-18.5</position>
<input>
<ID>IN_0</ID>379 </input>
<input>
<ID>IN_1</ID>381 </input>
<input>
<ID>IN_2</ID>380 </input>
<input>
<ID>IN_3</ID>378 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>223</ID>
<type>AA_REGISTER4</type>
<position>276,-1.5</position>
<output>
<ID>OUT_0</ID>379 </output>
<output>
<ID>OUT_1</ID>381 </output>
<output>
<ID>OUT_2</ID>380 </output>
<output>
<ID>OUT_3</ID>378 </output>
<input>
<ID>clear</ID>386 </input>
<input>
<ID>clock</ID>377 </input>
<input>
<ID>count_enable</ID>377 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>224</ID>
<type>AA_AND2</type>
<position>277,-9</position>
<input>
<ID>IN_0</ID>378 </input>
<input>
<ID>IN_1</ID>379 </input>
<output>
<ID>OUT</ID>386 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>225</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>274,-18.5</position>
<input>
<ID>IN_0</ID>383 </input>
<input>
<ID>IN_1</ID>385 </input>
<input>
<ID>IN_2</ID>384 </input>
<input>
<ID>IN_3</ID>382 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>226</ID>
<type>AA_REGISTER4</type>
<position>265.5,-1.5</position>
<output>
<ID>OUT_0</ID>383 </output>
<output>
<ID>OUT_1</ID>385 </output>
<output>
<ID>OUT_2</ID>384 </output>
<output>
<ID>OUT_3</ID>382 </output>
<input>
<ID>clear</ID>392 </input>
<input>
<ID>clock</ID>386 </input>
<input>
<ID>count_enable</ID>386 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>227</ID>
<type>AA_AND2</type>
<position>266.5,-9</position>
<input>
<ID>IN_0</ID>382 </input>
<input>
<ID>IN_1</ID>383 </input>
<output>
<ID>OUT</ID>392 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>228</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>263.5,-18.5</position>
<input>
<ID>IN_0</ID>388 </input>
<input>
<ID>IN_1</ID>390 </input>
<input>
<ID>IN_2</ID>389 </input>
<input>
<ID>IN_3</ID>387 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>229</ID>
<type>AA_REGISTER4</type>
<position>255,-1.5</position>
<output>
<ID>OUT_0</ID>388 </output>
<output>
<ID>OUT_1</ID>390 </output>
<output>
<ID>OUT_2</ID>389 </output>
<output>
<ID>OUT_3</ID>387 </output>
<input>
<ID>clear</ID>420 </input>
<input>
<ID>clock</ID>392 </input>
<input>
<ID>count_enable</ID>392 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>230</ID>
<type>AA_AND2</type>
<position>256,-9</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>388 </input>
<output>
<ID>OUT</ID>420 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>231</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>253,-18.5</position>
<input>
<ID>IN_0</ID>395 </input>
<input>
<ID>IN_1</ID>397 </input>
<input>
<ID>IN_2</ID>396 </input>
<input>
<ID>IN_3</ID>394 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>232</ID>
<type>AA_REGISTER4</type>
<position>244.5,-1.5</position>
<output>
<ID>OUT_0</ID>395 </output>
<output>
<ID>OUT_1</ID>397 </output>
<output>
<ID>OUT_2</ID>396 </output>
<output>
<ID>OUT_3</ID>394 </output>
<input>
<ID>clear</ID>421 </input>
<input>
<ID>clock</ID>420 </input>
<input>
<ID>count_enable</ID>420 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>233</ID>
<type>AA_AND2</type>
<position>245.5,-9</position>
<input>
<ID>IN_0</ID>394 </input>
<input>
<ID>IN_1</ID>395 </input>
<output>
<ID>OUT</ID>421 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>234</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>242.5,-18.5</position>
<input>
<ID>IN_0</ID>400 </input>
<input>
<ID>IN_1</ID>402 </input>
<input>
<ID>IN_2</ID>401 </input>
<input>
<ID>IN_3</ID>399 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>235</ID>
<type>AA_REGISTER4</type>
<position>234,-1.5</position>
<output>
<ID>OUT_0</ID>400 </output>
<output>
<ID>OUT_1</ID>402 </output>
<output>
<ID>OUT_2</ID>401 </output>
<output>
<ID>OUT_3</ID>399 </output>
<input>
<ID>clear</ID>403 </input>
<input>
<ID>clock</ID>421 </input>
<input>
<ID>count_enable</ID>421 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_AND2</type>
<position>235,-9</position>
<input>
<ID>IN_0</ID>399 </input>
<input>
<ID>IN_1</ID>400 </input>
<output>
<ID>OUT</ID>403 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>237</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>232,-18.5</position>
<input>
<ID>IN_0</ID>405 </input>
<input>
<ID>IN_1</ID>407 </input>
<input>
<ID>IN_2</ID>406 </input>
<input>
<ID>IN_3</ID>404 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>238</ID>
<type>AA_REGISTER4</type>
<position>223.5,-1.5</position>
<output>
<ID>OUT_0</ID>405 </output>
<output>
<ID>OUT_1</ID>407 </output>
<output>
<ID>OUT_2</ID>406 </output>
<output>
<ID>OUT_3</ID>404 </output>
<input>
<ID>clear</ID>412 </input>
<input>
<ID>clock</ID>403 </input>
<input>
<ID>count_enable</ID>403 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>239</ID>
<type>AA_AND2</type>
<position>224.5,-9</position>
<input>
<ID>IN_0</ID>404 </input>
<input>
<ID>IN_1</ID>405 </input>
<output>
<ID>OUT</ID>412 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>221.5,-18.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>411 </input>
<input>
<ID>IN_2</ID>410 </input>
<input>
<ID>IN_3</ID>408 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>241</ID>
<type>AA_REGISTER4</type>
<position>213,-1.5</position>
<output>
<ID>OUT_0</ID>409 </output>
<output>
<ID>OUT_1</ID>411 </output>
<output>
<ID>OUT_2</ID>410 </output>
<output>
<ID>OUT_3</ID>408 </output>
<input>
<ID>clear</ID>418 </input>
<input>
<ID>clock</ID>412 </input>
<input>
<ID>count_enable</ID>412 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>242</ID>
<type>AA_AND2</type>
<position>214,-9</position>
<input>
<ID>IN_0</ID>408 </input>
<input>
<ID>IN_1</ID>409 </input>
<output>
<ID>OUT</ID>418 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>243</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>211,-18.5</position>
<input>
<ID>IN_0</ID>414 </input>
<input>
<ID>IN_1</ID>416 </input>
<input>
<ID>IN_2</ID>415 </input>
<input>
<ID>IN_3</ID>413 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>244</ID>
<type>AA_REGISTER4</type>
<position>202.5,-1.5</position>
<output>
<ID>OUT_0</ID>414 </output>
<output>
<ID>OUT_1</ID>416 </output>
<output>
<ID>OUT_2</ID>415 </output>
<output>
<ID>OUT_3</ID>413 </output>
<input>
<ID>clear</ID>417 </input>
<input>
<ID>clock</ID>418 </input>
<input>
<ID>count_enable</ID>418 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>245</ID>
<type>AA_AND2</type>
<position>203.5,-9</position>
<input>
<ID>IN_0</ID>413 </input>
<input>
<ID>IN_1</ID>414 </input>
<output>
<ID>OUT</ID>417 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>246</ID>
<type>AA_REGISTER4</type>
<position>265.5,-28</position>
<output>
<ID>OUT_0</ID>356 </output>
<output>
<ID>OUT_1</ID>358 </output>
<output>
<ID>OUT_2</ID>357 </output>
<output>
<ID>OUT_3</ID>355 </output>
<input>
<ID>clear</ID>364 </input>
<input>
<ID>clock</ID>359 </input>
<input>
<ID>count_enable</ID>359 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>247</ID>
<type>AA_AND2</type>
<position>266.5,-35.5</position>
<input>
<ID>IN_0</ID>355 </input>
<input>
<ID>IN_1</ID>356 </input>
<output>
<ID>OUT</ID>364 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>248</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>263.5,-45</position>
<input>
<ID>IN_0</ID>361 </input>
<input>
<ID>IN_1</ID>363 </input>
<input>
<ID>IN_2</ID>362 </input>
<input>
<ID>IN_3</ID>360 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>249</ID>
<type>AA_REGISTER4</type>
<position>255,-28</position>
<output>
<ID>OUT_0</ID>361 </output>
<output>
<ID>OUT_1</ID>363 </output>
<output>
<ID>OUT_2</ID>362 </output>
<output>
<ID>OUT_3</ID>360 </output>
<input>
<ID>clear</ID>440 </input>
<input>
<ID>clock</ID>364 </input>
<input>
<ID>count_enable</ID>364 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_AND2</type>
<position>256,-35.5</position>
<input>
<ID>IN_0</ID>360 </input>
<input>
<ID>IN_1</ID>361 </input>
<output>
<ID>OUT</ID>440 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>251</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>253,-45</position>
<input>
<ID>IN_0</ID>372 </input>
<input>
<ID>IN_1</ID>398 </input>
<input>
<ID>IN_2</ID>391 </input>
<input>
<ID>IN_3</ID>366 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>252</ID>
<type>AA_REGISTER4</type>
<position>244.5,-28</position>
<output>
<ID>OUT_0</ID>372 </output>
<output>
<ID>OUT_1</ID>398 </output>
<output>
<ID>OUT_2</ID>391 </output>
<output>
<ID>OUT_3</ID>366 </output>
<input>
<ID>clear</ID>441 </input>
<input>
<ID>clock</ID>440 </input>
<input>
<ID>count_enable</ID>440 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_AND2</type>
<position>245.5,-35.5</position>
<input>
<ID>IN_0</ID>366 </input>
<input>
<ID>IN_1</ID>372 </input>
<output>
<ID>OUT</ID>441 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>254</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>242.5,-45</position>
<input>
<ID>IN_0</ID>422 </input>
<input>
<ID>IN_1</ID>424 </input>
<input>
<ID>IN_2</ID>423 </input>
<input>
<ID>IN_3</ID>419 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>255</ID>
<type>AA_REGISTER4</type>
<position>234,-28</position>
<output>
<ID>OUT_0</ID>422 </output>
<output>
<ID>OUT_1</ID>424 </output>
<output>
<ID>OUT_2</ID>423 </output>
<output>
<ID>OUT_3</ID>419 </output>
<input>
<ID>clear</ID>425 </input>
<input>
<ID>clock</ID>441 </input>
<input>
<ID>count_enable</ID>441 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>256</ID>
<type>AA_AND2</type>
<position>235,-35.5</position>
<input>
<ID>IN_0</ID>419 </input>
<input>
<ID>IN_1</ID>422 </input>
<output>
<ID>OUT</ID>425 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>257</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>232,-45</position>
<input>
<ID>IN_0</ID>427 </input>
<input>
<ID>IN_1</ID>429 </input>
<input>
<ID>IN_2</ID>428 </input>
<input>
<ID>IN_3</ID>426 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>258</ID>
<type>AA_REGISTER4</type>
<position>223.5,-28</position>
<output>
<ID>OUT_0</ID>427 </output>
<output>
<ID>OUT_1</ID>429 </output>
<output>
<ID>OUT_2</ID>428 </output>
<output>
<ID>OUT_3</ID>426 </output>
<input>
<ID>clear</ID>434 </input>
<input>
<ID>clock</ID>425 </input>
<input>
<ID>count_enable</ID>425 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>259</ID>
<type>AA_AND2</type>
<position>224.5,-35.5</position>
<input>
<ID>IN_0</ID>426 </input>
<input>
<ID>IN_1</ID>427 </input>
<output>
<ID>OUT</ID>434 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>260</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>221.5,-45</position>
<input>
<ID>IN_0</ID>431 </input>
<input>
<ID>IN_1</ID>433 </input>
<input>
<ID>IN_2</ID>432 </input>
<input>
<ID>IN_3</ID>430 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>261</ID>
<type>AA_REGISTER4</type>
<position>213,-28</position>
<output>
<ID>OUT_0</ID>431 </output>
<output>
<ID>OUT_1</ID>433 </output>
<output>
<ID>OUT_2</ID>432 </output>
<output>
<ID>OUT_3</ID>430 </output>
<input>
<ID>clear</ID>439 </input>
<input>
<ID>clock</ID>434 </input>
<input>
<ID>count_enable</ID>434 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>262</ID>
<type>AA_AND2</type>
<position>214,-35.5</position>
<input>
<ID>IN_0</ID>430 </input>
<input>
<ID>IN_1</ID>431 </input>
<output>
<ID>OUT</ID>439 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>263</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>211,-45</position>
<input>
<ID>IN_0</ID>436 </input>
<input>
<ID>IN_1</ID>438 </input>
<input>
<ID>IN_2</ID>437 </input>
<input>
<ID>IN_3</ID>435 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_REGISTER4</type>
<position>202.5,-28</position>
<output>
<ID>OUT_0</ID>436 </output>
<output>
<ID>OUT_1</ID>438 </output>
<output>
<ID>OUT_2</ID>437 </output>
<output>
<ID>OUT_3</ID>435 </output>
<input>
<ID>clear</ID>393 </input>
<input>
<ID>clock</ID>439 </input>
<input>
<ID>count_enable</ID>439 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_AND2</type>
<position>203.5,-35.5</position>
<input>
<ID>IN_0</ID>435 </input>
<input>
<ID>IN_1</ID>436 </input>
<output>
<ID>OUT</ID>393 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>266</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>305.5,8.5</position>
<input>
<ID>IN_0</ID>443 </input>
<input>
<ID>IN_1</ID>445 </input>
<input>
<ID>IN_2</ID>444 </input>
<input>
<ID>IN_3</ID>442 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>267</ID>
<type>AA_REGISTER4</type>
<position>297,25.5</position>
<output>
<ID>OUT_0</ID>443 </output>
<output>
<ID>OUT_1</ID>445 </output>
<output>
<ID>OUT_2</ID>444 </output>
<output>
<ID>OUT_3</ID>442 </output>
<input>
<ID>clear</ID>446 </input>
<input>
<ID>clock</ID>417 </input>
<input>
<ID>count_enable</ID>417 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>268</ID>
<type>AA_AND2</type>
<position>298,18</position>
<input>
<ID>IN_0</ID>442 </input>
<input>
<ID>IN_1</ID>443 </input>
<output>
<ID>OUT</ID>446 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>269</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>295,8.5</position>
<input>
<ID>IN_0</ID>448 </input>
<input>
<ID>IN_1</ID>450 </input>
<input>
<ID>IN_2</ID>449 </input>
<input>
<ID>IN_3</ID>447 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>270</ID>
<type>AA_REGISTER4</type>
<position>286.5,25.5</position>
<output>
<ID>OUT_0</ID>448 </output>
<output>
<ID>OUT_1</ID>450 </output>
<output>
<ID>OUT_2</ID>449 </output>
<output>
<ID>OUT_3</ID>447 </output>
<input>
<ID>clear</ID>451 </input>
<input>
<ID>clock</ID>446 </input>
<input>
<ID>count_enable</ID>446 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>271</ID>
<type>AA_AND2</type>
<position>287.5,18</position>
<input>
<ID>IN_0</ID>447 </input>
<input>
<ID>IN_1</ID>448 </input>
<output>
<ID>OUT</ID>451 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>272</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>284.5,8.5</position>
<input>
<ID>IN_0</ID>453 </input>
<input>
<ID>IN_1</ID>455 </input>
<input>
<ID>IN_2</ID>454 </input>
<input>
<ID>IN_3</ID>452 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>273</ID>
<type>AA_REGISTER4</type>
<position>276,25.5</position>
<output>
<ID>OUT_0</ID>453 </output>
<output>
<ID>OUT_1</ID>455 </output>
<output>
<ID>OUT_2</ID>454 </output>
<output>
<ID>OUT_3</ID>452 </output>
<input>
<ID>clear</ID>460 </input>
<input>
<ID>clock</ID>451 </input>
<input>
<ID>count_enable</ID>451 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>274</ID>
<type>AA_AND2</type>
<position>277,18</position>
<input>
<ID>IN_0</ID>452 </input>
<input>
<ID>IN_1</ID>453 </input>
<output>
<ID>OUT</ID>460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>275</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>274,8.5</position>
<input>
<ID>IN_0</ID>457 </input>
<input>
<ID>IN_1</ID>459 </input>
<input>
<ID>IN_2</ID>458 </input>
<input>
<ID>IN_3</ID>456 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>276</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>305.5,35</position>
<input>
<ID>IN_0</ID>469 </input>
<input>
<ID>IN_1</ID>471 </input>
<input>
<ID>IN_2</ID>470 </input>
<input>
<ID>IN_3</ID>468 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>277</ID>
<type>AA_REGISTER4</type>
<position>297,52</position>
<output>
<ID>OUT_0</ID>469 </output>
<output>
<ID>OUT_1</ID>471 </output>
<output>
<ID>OUT_2</ID>470 </output>
<output>
<ID>OUT_3</ID>468 </output>
<input>
<ID>clear</ID>472 </input>
<input>
<ID>clock</ID>494 </input>
<input>
<ID>count_enable</ID>494 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>278</ID>
<type>AA_AND2</type>
<position>298,44.5</position>
<input>
<ID>IN_0</ID>468 </input>
<input>
<ID>IN_1</ID>469 </input>
<output>
<ID>OUT</ID>472 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>279</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>295,35</position>
<input>
<ID>IN_0</ID>475 </input>
<input>
<ID>IN_1</ID>477 </input>
<input>
<ID>IN_2</ID>476 </input>
<input>
<ID>IN_3</ID>474 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>280</ID>
<type>AA_REGISTER4</type>
<position>286.5,52</position>
<output>
<ID>OUT_0</ID>475 </output>
<output>
<ID>OUT_1</ID>477 </output>
<output>
<ID>OUT_2</ID>476 </output>
<output>
<ID>OUT_3</ID>474 </output>
<input>
<ID>clear</ID>478 </input>
<input>
<ID>clock</ID>472 </input>
<input>
<ID>count_enable</ID>472 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>281</ID>
<type>AA_AND2</type>
<position>287.5,44.5</position>
<input>
<ID>IN_0</ID>474 </input>
<input>
<ID>IN_1</ID>475 </input>
<output>
<ID>OUT</ID>478 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>282</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>284.5,35</position>
<input>
<ID>IN_0</ID>480 </input>
<input>
<ID>IN_1</ID>482 </input>
<input>
<ID>IN_2</ID>481 </input>
<input>
<ID>IN_3</ID>479 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>283</ID>
<type>AA_REGISTER4</type>
<position>276,52</position>
<output>
<ID>OUT_0</ID>480 </output>
<output>
<ID>OUT_1</ID>482 </output>
<output>
<ID>OUT_2</ID>481 </output>
<output>
<ID>OUT_3</ID>479 </output>
<input>
<ID>clear</ID>487 </input>
<input>
<ID>clock</ID>478 </input>
<input>
<ID>count_enable</ID>478 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>284</ID>
<type>AA_AND2</type>
<position>277,44.5</position>
<input>
<ID>IN_0</ID>479 </input>
<input>
<ID>IN_1</ID>480 </input>
<output>
<ID>OUT</ID>487 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>285</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>274,35</position>
<input>
<ID>IN_0</ID>484 </input>
<input>
<ID>IN_1</ID>486 </input>
<input>
<ID>IN_2</ID>485 </input>
<input>
<ID>IN_3</ID>483 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>286</ID>
<type>AA_REGISTER4</type>
<position>265.5,52</position>
<output>
<ID>OUT_0</ID>484 </output>
<output>
<ID>OUT_1</ID>486 </output>
<output>
<ID>OUT_2</ID>485 </output>
<output>
<ID>OUT_3</ID>483 </output>
<input>
<ID>clear</ID>493 </input>
<input>
<ID>clock</ID>487 </input>
<input>
<ID>count_enable</ID>487 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>287</ID>
<type>AA_AND2</type>
<position>266.5,44.5</position>
<input>
<ID>IN_0</ID>483 </input>
<input>
<ID>IN_1</ID>484 </input>
<output>
<ID>OUT</ID>493 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>288</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>263.5,35</position>
<input>
<ID>IN_0</ID>489 </input>
<input>
<ID>IN_1</ID>491 </input>
<input>
<ID>IN_2</ID>490 </input>
<input>
<ID>IN_3</ID>488 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>289</ID>
<type>AA_REGISTER4</type>
<position>255,52</position>
<output>
<ID>OUT_0</ID>489 </output>
<output>
<ID>OUT_1</ID>491 </output>
<output>
<ID>OUT_2</ID>490 </output>
<output>
<ID>OUT_3</ID>488 </output>
<input>
<ID>clear</ID>521 </input>
<input>
<ID>clock</ID>493 </input>
<input>
<ID>count_enable</ID>493 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>290</ID>
<type>AA_AND2</type>
<position>256,44.5</position>
<input>
<ID>IN_0</ID>488 </input>
<input>
<ID>IN_1</ID>489 </input>
<output>
<ID>OUT</ID>521 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>291</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>253,35</position>
<input>
<ID>IN_0</ID>496 </input>
<input>
<ID>IN_1</ID>498 </input>
<input>
<ID>IN_2</ID>497 </input>
<input>
<ID>IN_3</ID>495 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>292</ID>
<type>AA_REGISTER4</type>
<position>244.5,52</position>
<output>
<ID>OUT_0</ID>496 </output>
<output>
<ID>OUT_1</ID>498 </output>
<output>
<ID>OUT_2</ID>497 </output>
<output>
<ID>OUT_3</ID>495 </output>
<input>
<ID>clear</ID>522 </input>
<input>
<ID>clock</ID>521 </input>
<input>
<ID>count_enable</ID>521 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>293</ID>
<type>AA_AND2</type>
<position>245.5,44.5</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>496 </input>
<output>
<ID>OUT</ID>522 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>294</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>242.5,35</position>
<input>
<ID>IN_0</ID>501 </input>
<input>
<ID>IN_1</ID>503 </input>
<input>
<ID>IN_2</ID>502 </input>
<input>
<ID>IN_3</ID>500 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>295</ID>
<type>AA_REGISTER4</type>
<position>234,52</position>
<output>
<ID>OUT_0</ID>501 </output>
<output>
<ID>OUT_1</ID>503 </output>
<output>
<ID>OUT_2</ID>502 </output>
<output>
<ID>OUT_3</ID>500 </output>
<input>
<ID>clear</ID>504 </input>
<input>
<ID>clock</ID>522 </input>
<input>
<ID>count_enable</ID>522 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>296</ID>
<type>AA_AND2</type>
<position>235,44.5</position>
<input>
<ID>IN_0</ID>500 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>504 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>297</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>232,35</position>
<input>
<ID>IN_0</ID>506 </input>
<input>
<ID>IN_1</ID>508 </input>
<input>
<ID>IN_2</ID>507 </input>
<input>
<ID>IN_3</ID>505 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>298</ID>
<type>AA_REGISTER4</type>
<position>223.5,52</position>
<output>
<ID>OUT_0</ID>506 </output>
<output>
<ID>OUT_1</ID>508 </output>
<output>
<ID>OUT_2</ID>507 </output>
<output>
<ID>OUT_3</ID>505 </output>
<input>
<ID>clear</ID>513 </input>
<input>
<ID>clock</ID>504 </input>
<input>
<ID>count_enable</ID>504 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>299</ID>
<type>AA_AND2</type>
<position>224.5,44.5</position>
<input>
<ID>IN_0</ID>505 </input>
<input>
<ID>IN_1</ID>506 </input>
<output>
<ID>OUT</ID>513 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>300</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>221.5,35</position>
<input>
<ID>IN_0</ID>510 </input>
<input>
<ID>IN_1</ID>512 </input>
<input>
<ID>IN_2</ID>511 </input>
<input>
<ID>IN_3</ID>509 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>301</ID>
<type>AA_REGISTER4</type>
<position>213,52</position>
<output>
<ID>OUT_0</ID>510 </output>
<output>
<ID>OUT_1</ID>512 </output>
<output>
<ID>OUT_2</ID>511 </output>
<output>
<ID>OUT_3</ID>509 </output>
<input>
<ID>clear</ID>519 </input>
<input>
<ID>clock</ID>513 </input>
<input>
<ID>count_enable</ID>513 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>302</ID>
<type>AA_AND2</type>
<position>214,44.5</position>
<input>
<ID>IN_0</ID>509 </input>
<input>
<ID>IN_1</ID>510 </input>
<output>
<ID>OUT</ID>519 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>303</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>211,35</position>
<input>
<ID>IN_0</ID>515 </input>
<input>
<ID>IN_1</ID>517 </input>
<input>
<ID>IN_2</ID>516 </input>
<input>
<ID>IN_3</ID>514 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>304</ID>
<type>AA_REGISTER4</type>
<position>202.5,52</position>
<output>
<ID>OUT_0</ID>515 </output>
<output>
<ID>OUT_1</ID>517 </output>
<output>
<ID>OUT_2</ID>516 </output>
<output>
<ID>OUT_3</ID>514 </output>
<input>
<ID>clear</ID>518 </input>
<input>
<ID>clock</ID>519 </input>
<input>
<ID>count_enable</ID>519 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>305</ID>
<type>AA_AND2</type>
<position>203.5,44.5</position>
<input>
<ID>IN_0</ID>514 </input>
<input>
<ID>IN_1</ID>515 </input>
<output>
<ID>OUT</ID>518 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>306</ID>
<type>AA_REGISTER4</type>
<position>265.5,25.5</position>
<output>
<ID>OUT_0</ID>457 </output>
<output>
<ID>OUT_1</ID>459 </output>
<output>
<ID>OUT_2</ID>458 </output>
<output>
<ID>OUT_3</ID>456 </output>
<input>
<ID>clear</ID>465 </input>
<input>
<ID>clock</ID>460 </input>
<input>
<ID>count_enable</ID>460 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>307</ID>
<type>AA_AND2</type>
<position>266.5,18</position>
<input>
<ID>IN_0</ID>456 </input>
<input>
<ID>IN_1</ID>457 </input>
<output>
<ID>OUT</ID>465 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>308</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>263.5,8.5</position>
<input>
<ID>IN_0</ID>462 </input>
<input>
<ID>IN_1</ID>464 </input>
<input>
<ID>IN_2</ID>463 </input>
<input>
<ID>IN_3</ID>461 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>309</ID>
<type>AA_REGISTER4</type>
<position>255,25.5</position>
<output>
<ID>OUT_0</ID>462 </output>
<output>
<ID>OUT_1</ID>464 </output>
<output>
<ID>OUT_2</ID>463 </output>
<output>
<ID>OUT_3</ID>461 </output>
<input>
<ID>clear</ID>541 </input>
<input>
<ID>clock</ID>465 </input>
<input>
<ID>count_enable</ID>465 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>310</ID>
<type>AA_AND2</type>
<position>256,18</position>
<input>
<ID>IN_0</ID>461 </input>
<input>
<ID>IN_1</ID>462 </input>
<output>
<ID>OUT</ID>541 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>311</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>253,8.5</position>
<input>
<ID>IN_0</ID>473 </input>
<input>
<ID>IN_1</ID>499 </input>
<input>
<ID>IN_2</ID>492 </input>
<input>
<ID>IN_3</ID>467 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>312</ID>
<type>AA_REGISTER4</type>
<position>244.5,25.5</position>
<output>
<ID>OUT_0</ID>473 </output>
<output>
<ID>OUT_1</ID>499 </output>
<output>
<ID>OUT_2</ID>492 </output>
<output>
<ID>OUT_3</ID>467 </output>
<input>
<ID>clear</ID>542 </input>
<input>
<ID>clock</ID>541 </input>
<input>
<ID>count_enable</ID>541 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>313</ID>
<type>AA_AND2</type>
<position>245.5,18</position>
<input>
<ID>IN_0</ID>467 </input>
<input>
<ID>IN_1</ID>473 </input>
<output>
<ID>OUT</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>314</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>242.5,8.5</position>
<input>
<ID>IN_0</ID>523 </input>
<input>
<ID>IN_1</ID>525 </input>
<input>
<ID>IN_2</ID>524 </input>
<input>
<ID>IN_3</ID>520 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>315</ID>
<type>AA_REGISTER4</type>
<position>234,25.5</position>
<output>
<ID>OUT_0</ID>523 </output>
<output>
<ID>OUT_1</ID>525 </output>
<output>
<ID>OUT_2</ID>524 </output>
<output>
<ID>OUT_3</ID>520 </output>
<input>
<ID>clear</ID>526 </input>
<input>
<ID>clock</ID>542 </input>
<input>
<ID>count_enable</ID>542 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>316</ID>
<type>AA_AND2</type>
<position>235,18</position>
<input>
<ID>IN_0</ID>520 </input>
<input>
<ID>IN_1</ID>523 </input>
<output>
<ID>OUT</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>317</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>232,8.5</position>
<input>
<ID>IN_0</ID>528 </input>
<input>
<ID>IN_1</ID>530 </input>
<input>
<ID>IN_2</ID>529 </input>
<input>
<ID>IN_3</ID>527 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>318</ID>
<type>AA_REGISTER4</type>
<position>223.5,25.5</position>
<output>
<ID>OUT_0</ID>528 </output>
<output>
<ID>OUT_1</ID>530 </output>
<output>
<ID>OUT_2</ID>529 </output>
<output>
<ID>OUT_3</ID>527 </output>
<input>
<ID>clear</ID>535 </input>
<input>
<ID>clock</ID>526 </input>
<input>
<ID>count_enable</ID>526 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>319</ID>
<type>AA_AND2</type>
<position>224.5,18</position>
<input>
<ID>IN_0</ID>527 </input>
<input>
<ID>IN_1</ID>528 </input>
<output>
<ID>OUT</ID>535 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>320</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>221.5,8.5</position>
<input>
<ID>IN_0</ID>532 </input>
<input>
<ID>IN_1</ID>534 </input>
<input>
<ID>IN_2</ID>533 </input>
<input>
<ID>IN_3</ID>531 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>321</ID>
<type>AA_REGISTER4</type>
<position>213,25.5</position>
<output>
<ID>OUT_0</ID>532 </output>
<output>
<ID>OUT_1</ID>534 </output>
<output>
<ID>OUT_2</ID>533 </output>
<output>
<ID>OUT_3</ID>531 </output>
<input>
<ID>clear</ID>540 </input>
<input>
<ID>clock</ID>535 </input>
<input>
<ID>count_enable</ID>535 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>322</ID>
<type>AA_AND2</type>
<position>214,18</position>
<input>
<ID>IN_0</ID>531 </input>
<input>
<ID>IN_1</ID>532 </input>
<output>
<ID>OUT</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>323</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>211,8.5</position>
<input>
<ID>IN_0</ID>537 </input>
<input>
<ID>IN_1</ID>539 </input>
<input>
<ID>IN_2</ID>538 </input>
<input>
<ID>IN_3</ID>536 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>324</ID>
<type>AA_REGISTER4</type>
<position>202.5,25.5</position>
<output>
<ID>OUT_0</ID>537 </output>
<output>
<ID>OUT_1</ID>539 </output>
<output>
<ID>OUT_2</ID>538 </output>
<output>
<ID>OUT_3</ID>536 </output>
<input>
<ID>clear</ID>494 </input>
<input>
<ID>clock</ID>540 </input>
<input>
<ID>count_enable</ID>540 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>325</ID>
<type>AA_AND2</type>
<position>203.5,18</position>
<input>
<ID>IN_0</ID>536 </input>
<input>
<ID>IN_1</ID>537 </input>
<output>
<ID>OUT</ID>494 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,-205,303.5,-188</points>
<connection>
<GID>5</GID>
<name>IN_3</name></connection>
<intersection>-201 1</intersection>
<intersection>-188 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>298,-201,303.5,-201</points>
<intersection>298 17</intersection>
<intersection>303.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>302,-188,303.5,-188</points>
<connection>
<GID>7</GID>
<name>OUT_3</name></connection>
<intersection>303.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>298,-201,298,-200.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>-201 1</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-208,302,-191</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-208 5</intersection>
<intersection>-200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>300,-200.5,302,-200.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>302 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>302,-208,303.5,-208</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>302 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303,-206,303,-189</points>
<intersection>-206 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303,-206,303.5,-206</points>
<connection>
<GID>5</GID>
<name>IN_2</name></connection>
<intersection>303 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>302,-189,303,-189</points>
<connection>
<GID>7</GID>
<name>OUT_2</name></connection>
<intersection>303 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,-207,302.5,-190</points>
<intersection>-207 3</intersection>
<intersection>-190 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>302,-190,302.5,-190</points>
<connection>
<GID>7</GID>
<name>OUT_1</name></connection>
<intersection>302.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>302.5,-207,303.5,-207</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>302.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>299,-194.5,299,-194</points>
<connection>
<GID>7</GID>
<name>clear</name></connection>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>-194.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>283,-194.5,299,-194.5</points>
<intersection>283 2</intersection>
<intersection>286.5 7</intersection>
<intersection>299 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>283,-194.5,283,-184.5</points>
<intersection>-194.5 1</intersection>
<intersection>-184.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>283,-184.5,287.5,-184.5</points>
<intersection>283 2</intersection>
<intersection>287.5 10</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>286.5,-194.5,286.5,-194</points>
<connection>
<GID>30</GID>
<name>clock</name></connection>
<intersection>-194.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>287.5,-185,287.5,-184.5</points>
<connection>
<GID>30</GID>
<name>count_enable</name></connection>
<intersection>-184.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-205,293,-188</points>
<connection>
<GID>17</GID>
<name>IN_3</name></connection>
<intersection>-201 1</intersection>
<intersection>-188 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287.5,-201,293,-201</points>
<intersection>287.5 17</intersection>
<intersection>293 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>291.5,-188,293,-188</points>
<connection>
<GID>30</GID>
<name>OUT_3</name></connection>
<intersection>293 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>287.5,-201,287.5,-200.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-201 1</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,-208,291.5,-191</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>-208 5</intersection>
<intersection>-200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>289.5,-200.5,291.5,-200.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>291.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>291.5,-208,293,-208</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,-206,292.5,-189</points>
<intersection>-206 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>292.5,-206,293,-206</points>
<connection>
<GID>17</GID>
<name>IN_2</name></connection>
<intersection>292.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>291.5,-189,292.5,-189</points>
<connection>
<GID>30</GID>
<name>OUT_2</name></connection>
<intersection>292.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,-207,292,-190</points>
<intersection>-207 3</intersection>
<intersection>-190 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>291.5,-190,292,-190</points>
<connection>
<GID>30</GID>
<name>OUT_1</name></connection>
<intersection>292 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>292,-207,293,-207</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>292 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288.5,-194.5,288.5,-194</points>
<connection>
<GID>30</GID>
<name>clear</name></connection>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>-194.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>272.5,-194.5,288.5,-194.5</points>
<intersection>272.5 2</intersection>
<intersection>276 12</intersection>
<intersection>288.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>272.5,-194.5,272.5,-185</points>
<intersection>-194.5 1</intersection>
<intersection>-185 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>272.5,-185,277,-185</points>
<connection>
<GID>33</GID>
<name>count_enable</name></connection>
<intersection>272.5 2</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>276,-194.5,276,-194</points>
<connection>
<GID>33</GID>
<name>clock</name></connection>
<intersection>-194.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282.5,-205,282.5,-188</points>
<connection>
<GID>32</GID>
<name>IN_3</name></connection>
<intersection>-201 1</intersection>
<intersection>-188 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>277,-201,282.5,-201</points>
<intersection>277 17</intersection>
<intersection>282.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281,-188,282.5,-188</points>
<connection>
<GID>33</GID>
<name>OUT_3</name></connection>
<intersection>282.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>277,-201,277,-200.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>-201 1</intersection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,-208,281,-191</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>-208 5</intersection>
<intersection>-200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>279,-200.5,281,-200.5</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>281 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>281,-208,282.5,-208</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>281 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-206,282,-189</points>
<intersection>-206 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282,-206,282.5,-206</points>
<connection>
<GID>32</GID>
<name>IN_2</name></connection>
<intersection>282 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281,-189,282,-189</points>
<connection>
<GID>33</GID>
<name>OUT_2</name></connection>
<intersection>282 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-207,281.5,-190</points>
<intersection>-207 3</intersection>
<intersection>-190 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>281,-190,281.5,-190</points>
<connection>
<GID>33</GID>
<name>OUT_1</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>281.5,-207,282.5,-207</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272,-205,272,-188</points>
<connection>
<GID>35</GID>
<name>IN_3</name></connection>
<intersection>-201 1</intersection>
<intersection>-188 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266.5,-201,272,-201</points>
<intersection>266.5 17</intersection>
<intersection>272 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>270.5,-188,272,-188</points>
<connection>
<GID>66</GID>
<name>OUT_3</name></connection>
<intersection>272 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>266.5,-201,266.5,-200.5</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>-201 1</intersection></vsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-208,270.5,-191</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>-208 5</intersection>
<intersection>-200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>268.5,-200.5,270.5,-200.5</points>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>270.5,-208,272,-208</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,-206,271.5,-189</points>
<intersection>-206 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>271.5,-206,272,-206</points>
<connection>
<GID>35</GID>
<name>IN_2</name></connection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>270.5,-189,271.5,-189</points>
<connection>
<GID>66</GID>
<name>OUT_2</name></connection>
<intersection>271.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-207,271,-190</points>
<intersection>-207 3</intersection>
<intersection>-190 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>270.5,-190,271,-190</points>
<connection>
<GID>66</GID>
<name>OUT_1</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>271,-207,272,-207</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>271 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262,-194.5,262,-184.5</points>
<intersection>-194.5 4</intersection>
<intersection>-184.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>262,-184.5,266.5,-184.5</points>
<intersection>262 0</intersection>
<intersection>266.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>262,-194.5,278,-194.5</points>
<intersection>262 0</intersection>
<intersection>265.5 7</intersection>
<intersection>278 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>278,-194.5,278,-194</points>
<connection>
<GID>33</GID>
<name>clear</name></connection>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>-194.5 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>265.5,-194.5,265.5,-194</points>
<connection>
<GID>66</GID>
<name>clock</name></connection>
<intersection>-194.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>266.5,-185,266.5,-184.5</points>
<connection>
<GID>66</GID>
<name>count_enable</name></connection>
<intersection>-184.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,-205,261.5,-188</points>
<connection>
<GID>68</GID>
<name>IN_3</name></connection>
<intersection>-201 1</intersection>
<intersection>-188 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>256,-201,261.5,-201</points>
<intersection>256 17</intersection>
<intersection>261.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>260,-188,261.5,-188</points>
<connection>
<GID>69</GID>
<name>OUT_3</name></connection>
<intersection>261.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>256,-201,256,-200.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>-201 1</intersection></vsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-208,260,-191</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<intersection>-208 5</intersection>
<intersection>-200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>258,-200.5,260,-200.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>260,-208,261.5,-208</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,-206,261,-189</points>
<intersection>-206 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261,-206,261.5,-206</points>
<connection>
<GID>68</GID>
<name>IN_2</name></connection>
<intersection>261 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>260,-189,261,-189</points>
<connection>
<GID>69</GID>
<name>OUT_2</name></connection>
<intersection>261 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,-207,260.5,-190</points>
<intersection>-207 3</intersection>
<intersection>-190 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>260,-190,260.5,-190</points>
<connection>
<GID>69</GID>
<name>OUT_1</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>260.5,-207,261.5,-207</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>260.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251.5,-194,251.5,-184.5</points>
<intersection>-194 4</intersection>
<intersection>-184.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>251.5,-184.5,256,-184.5</points>
<intersection>251.5 0</intersection>
<intersection>256 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>251.5,-194,267.5,-194</points>
<connection>
<GID>69</GID>
<name>clock</name></connection>
<intersection>251.5 0</intersection>
<intersection>267.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>267.5,-194.5,267.5,-194</points>
<connection>
<GID>66</GID>
<name>clear</name></connection>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<intersection>-194 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>256,-185,256,-184.5</points>
<connection>
<GID>69</GID>
<name>count_enable</name></connection>
<intersection>-184.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293.5,-194,293.5,-184.5</points>
<intersection>-194 4</intersection>
<intersection>-184.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>293.5,-184.5,298,-184.5</points>
<intersection>293.5 0</intersection>
<intersection>298 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293.5,-194,297,-194</points>
<connection>
<GID>7</GID>
<name>clock</name></connection>
<intersection>293.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>298,-185,298,-184.5</points>
<connection>
<GID>7</GID>
<name>count_enable</name></connection>
<intersection>-184.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,-205,251,-188</points>
<connection>
<GID>71</GID>
<name>IN_3</name></connection>
<intersection>-201 1</intersection>
<intersection>-188 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245.5,-201,251,-201</points>
<intersection>245.5 17</intersection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>249.5,-188,251,-188</points>
<connection>
<GID>72</GID>
<name>OUT_3</name></connection>
<intersection>251 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>245.5,-201,245.5,-200.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>-201 1</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,-178.5,303.5,-161.5</points>
<connection>
<GID>36</GID>
<name>IN_3</name></connection>
<intersection>-174.5 1</intersection>
<intersection>-161.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>298,-174.5,303.5,-174.5</points>
<intersection>298 17</intersection>
<intersection>303.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>302,-161.5,303.5,-161.5</points>
<connection>
<GID>37</GID>
<name>OUT_3</name></connection>
<intersection>303.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>298,-174.5,298,-174</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>-174.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-181.5,302,-164.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>-181.5 5</intersection>
<intersection>-174 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>300,-174,302,-174</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>302 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>302,-181.5,303.5,-181.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>302 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303,-179.5,303,-162.5</points>
<intersection>-179.5 1</intersection>
<intersection>-162.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303,-179.5,303.5,-179.5</points>
<connection>
<GID>36</GID>
<name>IN_2</name></connection>
<intersection>303 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>302,-162.5,303,-162.5</points>
<connection>
<GID>37</GID>
<name>OUT_2</name></connection>
<intersection>303 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,-180.5,302.5,-163.5</points>
<intersection>-180.5 3</intersection>
<intersection>-163.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>302,-163.5,302.5,-163.5</points>
<connection>
<GID>37</GID>
<name>OUT_1</name></connection>
<intersection>302.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>302.5,-180.5,303.5,-180.5</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>302.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>299,-168,299,-167.5</points>
<connection>
<GID>37</GID>
<name>clear</name></connection>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>-168 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>283,-168,299,-168</points>
<intersection>283 2</intersection>
<intersection>286.5 7</intersection>
<intersection>299 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>283,-168,283,-158</points>
<intersection>-168 1</intersection>
<intersection>-158 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>283,-158,287.5,-158</points>
<intersection>283 2</intersection>
<intersection>287.5 10</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>286.5,-168,286.5,-167.5</points>
<connection>
<GID>40</GID>
<name>clock</name></connection>
<intersection>-168 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>287.5,-158.5,287.5,-158</points>
<connection>
<GID>40</GID>
<name>count_enable</name></connection>
<intersection>-158 5</intersection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,-208,249.5,-191</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>-208 5</intersection>
<intersection>-200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>247.5,-200.5,249.5,-200.5</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>249.5,-208,251,-208</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-178.5,293,-161.5</points>
<connection>
<GID>39</GID>
<name>IN_3</name></connection>
<intersection>-174.5 1</intersection>
<intersection>-161.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287.5,-174.5,293,-174.5</points>
<intersection>287.5 17</intersection>
<intersection>293 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>291.5,-161.5,293,-161.5</points>
<connection>
<GID>40</GID>
<name>OUT_3</name></connection>
<intersection>293 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>287.5,-174.5,287.5,-174</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>-174.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,-181.5,291.5,-164.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>-181.5 5</intersection>
<intersection>-174 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>289.5,-174,291.5,-174</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>291.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>291.5,-181.5,293,-181.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,-179.5,292.5,-162.5</points>
<intersection>-179.5 1</intersection>
<intersection>-162.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>292.5,-179.5,293,-179.5</points>
<connection>
<GID>39</GID>
<name>IN_2</name></connection>
<intersection>292.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>291.5,-162.5,292.5,-162.5</points>
<connection>
<GID>40</GID>
<name>OUT_2</name></connection>
<intersection>292.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,-180.5,292,-163.5</points>
<intersection>-180.5 3</intersection>
<intersection>-163.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>291.5,-163.5,292,-163.5</points>
<connection>
<GID>40</GID>
<name>OUT_1</name></connection>
<intersection>292 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>292,-180.5,293,-180.5</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>292 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288.5,-168,288.5,-167.5</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<connection>
<GID>40</GID>
<name>clear</name></connection>
<intersection>-167.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>272.5,-167.5,288.5,-167.5</points>
<connection>
<GID>43</GID>
<name>clock</name></connection>
<intersection>272.5 2</intersection>
<intersection>288.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>272.5,-167.5,272.5,-158</points>
<intersection>-167.5 1</intersection>
<intersection>-158 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>272.5,-158,277,-158</points>
<intersection>272.5 2</intersection>
<intersection>277 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>277,-158.5,277,-158</points>
<connection>
<GID>43</GID>
<name>count_enable</name></connection>
<intersection>-158 5</intersection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282.5,-178.5,282.5,-161.5</points>
<connection>
<GID>42</GID>
<name>IN_3</name></connection>
<intersection>-174.5 1</intersection>
<intersection>-161.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>277,-174.5,282.5,-174.5</points>
<intersection>277 17</intersection>
<intersection>282.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281,-161.5,282.5,-161.5</points>
<connection>
<GID>43</GID>
<name>OUT_3</name></connection>
<intersection>282.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>277,-174.5,277,-174</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-174.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,-181.5,281,-164.5</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>-181.5 5</intersection>
<intersection>-174 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>279,-174,281,-174</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>281 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>281,-181.5,282.5,-181.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>281 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-179.5,282,-162.5</points>
<intersection>-179.5 1</intersection>
<intersection>-162.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282,-179.5,282.5,-179.5</points>
<connection>
<GID>42</GID>
<name>IN_2</name></connection>
<intersection>282 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281,-162.5,282,-162.5</points>
<connection>
<GID>43</GID>
<name>OUT_2</name></connection>
<intersection>282 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-180.5,281.5,-163.5</points>
<intersection>-180.5 3</intersection>
<intersection>-163.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>281,-163.5,281.5,-163.5</points>
<connection>
<GID>43</GID>
<name>OUT_1</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>281.5,-180.5,282.5,-180.5</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272,-178.5,272,-161.5</points>
<connection>
<GID>45</GID>
<name>IN_3</name></connection>
<intersection>-174.5 1</intersection>
<intersection>-161.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266.5,-174.5,272,-174.5</points>
<intersection>266.5 17</intersection>
<intersection>272 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>270.5,-161.5,272,-161.5</points>
<connection>
<GID>46</GID>
<name>OUT_3</name></connection>
<intersection>272 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>266.5,-174.5,266.5,-174</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>-174.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-181.5,270.5,-164.5</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>-181.5 5</intersection>
<intersection>-174 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>268.5,-174,270.5,-174</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>270.5,-181.5,272,-181.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,-179.5,271.5,-162.5</points>
<intersection>-179.5 1</intersection>
<intersection>-162.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>271.5,-179.5,272,-179.5</points>
<connection>
<GID>45</GID>
<name>IN_2</name></connection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>270.5,-162.5,271.5,-162.5</points>
<connection>
<GID>46</GID>
<name>OUT_2</name></connection>
<intersection>271.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-180.5,271,-163.5</points>
<intersection>-180.5 3</intersection>
<intersection>-163.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>270.5,-163.5,271,-163.5</points>
<connection>
<GID>46</GID>
<name>OUT_1</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>271,-180.5,272,-180.5</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>271 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262,-168,262,-158</points>
<intersection>-168 4</intersection>
<intersection>-158 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>262,-158,266.5,-158</points>
<intersection>262 0</intersection>
<intersection>266.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>262,-168,278,-168</points>
<intersection>262 0</intersection>
<intersection>265.5 7</intersection>
<intersection>278 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>278,-168,278,-167.5</points>
<connection>
<GID>43</GID>
<name>clear</name></connection>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>-168 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>265.5,-168,265.5,-167.5</points>
<connection>
<GID>46</GID>
<name>clock</name></connection>
<intersection>-168 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>266.5,-158.5,266.5,-158</points>
<connection>
<GID>46</GID>
<name>count_enable</name></connection>
<intersection>-158 3</intersection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,-178.5,261.5,-161.5</points>
<connection>
<GID>48</GID>
<name>IN_3</name></connection>
<intersection>-174.5 1</intersection>
<intersection>-161.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>256,-174.5,261.5,-174.5</points>
<intersection>256 17</intersection>
<intersection>261.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>260,-161.5,261.5,-161.5</points>
<connection>
<GID>49</GID>
<name>OUT_3</name></connection>
<intersection>261.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>256,-174.5,256,-174</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>-174.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-181.5,260,-164.5</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>-181.5 5</intersection>
<intersection>-174 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>258,-174,260,-174</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>260,-181.5,261.5,-181.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,-179.5,261,-162.5</points>
<intersection>-179.5 1</intersection>
<intersection>-162.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261,-179.5,261.5,-179.5</points>
<connection>
<GID>48</GID>
<name>IN_2</name></connection>
<intersection>261 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>260,-162.5,261,-162.5</points>
<connection>
<GID>49</GID>
<name>OUT_2</name></connection>
<intersection>261 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,-180.5,260.5,-163.5</points>
<intersection>-180.5 3</intersection>
<intersection>-163.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>260,-163.5,260.5,-163.5</points>
<connection>
<GID>49</GID>
<name>OUT_1</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>260.5,-180.5,261.5,-180.5</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>260.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,-206,250.5,-189</points>
<intersection>-206 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250.5,-206,251,-206</points>
<connection>
<GID>71</GID>
<name>IN_2</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>249.5,-189,250.5,-189</points>
<connection>
<GID>72</GID>
<name>OUT_2</name></connection>
<intersection>250.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251.5,-167.5,251.5,-158</points>
<intersection>-167.5 4</intersection>
<intersection>-158 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>251.5,-158,256,-158</points>
<intersection>251.5 0</intersection>
<intersection>256 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>251.5,-167.5,267.5,-167.5</points>
<connection>
<GID>49</GID>
<name>clock</name></connection>
<intersection>251.5 0</intersection>
<intersection>267.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>267.5,-168,267.5,-167.5</points>
<connection>
<GID>46</GID>
<name>clear</name></connection>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>-167.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>256,-158.5,256,-158</points>
<connection>
<GID>49</GID>
<name>count_enable</name></connection>
<intersection>-158 3</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293.5,-167.5,293.5,-158</points>
<intersection>-167.5 4</intersection>
<intersection>-158 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>293.5,-158,298,-158</points>
<intersection>293.5 0</intersection>
<intersection>298 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293.5,-167.5,297,-167.5</points>
<connection>
<GID>37</GID>
<name>clock</name></connection>
<intersection>293.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>298,-158.5,298,-157</points>
<connection>
<GID>37</GID>
<name>count_enable</name></connection>
<intersection>-158 3</intersection>
<intersection>-157 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>197,-157,298,-157</points>
<intersection>197 7</intersection>
<intersection>298 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>197,-194.5,197,-157</points>
<intersection>-194.5 8</intersection>
<intersection>-157 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>197,-194.5,204.5,-194.5</points>
<connection>
<GID>85</GID>
<name>OUT</name></connection>
<intersection>197 7</intersection>
<intersection>204.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>204.5,-194.5,204.5,-194</points>
<connection>
<GID>84</GID>
<name>clear</name></connection>
<intersection>-194.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,-178.5,251,-161.5</points>
<connection>
<GID>51</GID>
<name>IN_3</name></connection>
<intersection>-174.5 1</intersection>
<intersection>-161.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245.5,-174.5,251,-174.5</points>
<intersection>245.5 17</intersection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>249.5,-161.5,251,-161.5</points>
<connection>
<GID>52</GID>
<name>OUT_3</name></connection>
<intersection>251 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>245.5,-174.5,245.5,-174</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>-174.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,-181.5,249.5,-164.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>-181.5 5</intersection>
<intersection>-174 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>247.5,-174,249.5,-174</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>249.5,-181.5,251,-181.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,-179.5,250.5,-162.5</points>
<intersection>-179.5 1</intersection>
<intersection>-162.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250.5,-179.5,251,-179.5</points>
<connection>
<GID>51</GID>
<name>IN_2</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>249.5,-162.5,250.5,-162.5</points>
<connection>
<GID>52</GID>
<name>OUT_2</name></connection>
<intersection>250.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,-180.5,250,-163.5</points>
<intersection>-180.5 3</intersection>
<intersection>-163.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>249.5,-163.5,250,-163.5</points>
<connection>
<GID>52</GID>
<name>OUT_1</name></connection>
<intersection>250 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>250,-180.5,251,-180.5</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>250 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,-207,250,-190</points>
<intersection>-207 3</intersection>
<intersection>-190 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>249.5,-190,250,-190</points>
<connection>
<GID>72</GID>
<name>OUT_1</name></connection>
<intersection>250 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>250,-207,251,-207</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<intersection>250 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240.5,-178.5,240.5,-161.5</points>
<connection>
<GID>54</GID>
<name>IN_3</name></connection>
<intersection>-174.5 1</intersection>
<intersection>-161.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235,-174.5,240.5,-174.5</points>
<intersection>235 17</intersection>
<intersection>240.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>239,-161.5,240.5,-161.5</points>
<connection>
<GID>55</GID>
<name>OUT_3</name></connection>
<intersection>240.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>235,-174.5,235,-174</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>-174.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,-181.5,239,-164.5</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>-181.5 5</intersection>
<intersection>-174 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>237,-174,239,-174</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>239 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>239,-181.5,240.5,-181.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>239 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-179.5,240,-162.5</points>
<intersection>-179.5 1</intersection>
<intersection>-162.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240,-179.5,240.5,-179.5</points>
<connection>
<GID>54</GID>
<name>IN_2</name></connection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>239,-162.5,240,-162.5</points>
<connection>
<GID>55</GID>
<name>OUT_2</name></connection>
<intersection>240 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239.5,-180.5,239.5,-163.5</points>
<intersection>-180.5 3</intersection>
<intersection>-163.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>239,-163.5,239.5,-163.5</points>
<connection>
<GID>55</GID>
<name>OUT_1</name></connection>
<intersection>239.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>239.5,-180.5,240.5,-180.5</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>239.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,-168,236,-167.5</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<connection>
<GID>55</GID>
<name>clear</name></connection>
<intersection>-168 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>220,-168,236,-168</points>
<intersection>220 2</intersection>
<intersection>223.5 10</intersection>
<intersection>236 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-168,220,-158</points>
<intersection>-168 1</intersection>
<intersection>-158 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>220,-158,224.5,-158</points>
<intersection>220 2</intersection>
<intersection>224.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>224.5,-158.5,224.5,-158</points>
<connection>
<GID>58</GID>
<name>count_enable</name></connection>
<intersection>-158 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>223.5,-168,223.5,-167.5</points>
<connection>
<GID>58</GID>
<name>clock</name></connection>
<intersection>-168 1</intersection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,-178.5,230,-161.5</points>
<connection>
<GID>57</GID>
<name>IN_3</name></connection>
<intersection>-174.5 1</intersection>
<intersection>-161.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>224.5,-174.5,230,-174.5</points>
<intersection>224.5 17</intersection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228.5,-161.5,230,-161.5</points>
<connection>
<GID>58</GID>
<name>OUT_3</name></connection>
<intersection>230 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>224.5,-174.5,224.5,-174</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>-174.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,-181.5,228.5,-164.5</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>-181.5 5</intersection>
<intersection>-174 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-174,228.5,-174</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>228.5,-181.5,230,-181.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>228.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,-179.5,229.5,-162.5</points>
<intersection>-179.5 1</intersection>
<intersection>-162.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229.5,-179.5,230,-179.5</points>
<connection>
<GID>57</GID>
<name>IN_2</name></connection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228.5,-162.5,229.5,-162.5</points>
<connection>
<GID>58</GID>
<name>OUT_2</name></connection>
<intersection>229.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-180.5,229,-163.5</points>
<intersection>-180.5 3</intersection>
<intersection>-163.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>228.5,-163.5,229,-163.5</points>
<connection>
<GID>58</GID>
<name>OUT_1</name></connection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>229,-180.5,230,-180.5</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>229 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,-178.5,219.5,-161.5</points>
<connection>
<GID>60</GID>
<name>IN_3</name></connection>
<intersection>-174.5 1</intersection>
<intersection>-161.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>214,-174.5,219.5,-174.5</points>
<intersection>214 17</intersection>
<intersection>219.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>218,-161.5,219.5,-161.5</points>
<connection>
<GID>61</GID>
<name>OUT_3</name></connection>
<intersection>219.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>214,-174.5,214,-174</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-174.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-181.5,218,-164.5</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<intersection>-181.5 5</intersection>
<intersection>-174 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-174,218,-174</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>218,-181.5,219.5,-181.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-179.5,219,-162.5</points>
<intersection>-179.5 1</intersection>
<intersection>-162.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,-179.5,219.5,-179.5</points>
<connection>
<GID>60</GID>
<name>IN_2</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>218,-162.5,219,-162.5</points>
<connection>
<GID>61</GID>
<name>OUT_2</name></connection>
<intersection>219 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-180.5,218.5,-163.5</points>
<intersection>-180.5 3</intersection>
<intersection>-163.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>218,-163.5,218.5,-163.5</points>
<connection>
<GID>61</GID>
<name>OUT_1</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>218.5,-180.5,219.5,-180.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>218.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209.5,-167.5,209.5,-158</points>
<intersection>-167.5 4</intersection>
<intersection>-158 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>209.5,-158,214,-158</points>
<intersection>209.5 0</intersection>
<intersection>214 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>209.5,-167.5,225.5,-167.5</points>
<connection>
<GID>61</GID>
<name>clock</name></connection>
<intersection>209.5 0</intersection>
<intersection>225.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>225.5,-168,225.5,-167.5</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<connection>
<GID>58</GID>
<name>clear</name></connection>
<intersection>-167.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>214,-158.5,214,-158</points>
<connection>
<GID>61</GID>
<name>count_enable</name></connection>
<intersection>-158 3</intersection></vsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209,-178.5,209,-161.5</points>
<connection>
<GID>63</GID>
<name>IN_3</name></connection>
<intersection>-174.5 1</intersection>
<intersection>-161.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203.5,-174.5,209,-174.5</points>
<intersection>203.5 17</intersection>
<intersection>209 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207.5,-161.5,209,-161.5</points>
<connection>
<GID>64</GID>
<name>OUT_3</name></connection>
<intersection>209 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>203.5,-174.5,203.5,-174</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>-174.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,-181.5,207.5,-164.5</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>-181.5 5</intersection>
<intersection>-174 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>205.5,-174,207.5,-174</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<intersection>207.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>207.5,-181.5,209,-181.5</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>207.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-179.5,208.5,-162.5</points>
<intersection>-179.5 1</intersection>
<intersection>-162.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208.5,-179.5,209,-179.5</points>
<connection>
<GID>63</GID>
<name>IN_2</name></connection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207.5,-162.5,208.5,-162.5</points>
<connection>
<GID>64</GID>
<name>OUT_2</name></connection>
<intersection>208.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-180.5,208,-163.5</points>
<intersection>-180.5 3</intersection>
<intersection>-163.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>207.5,-163.5,208,-163.5</points>
<connection>
<GID>64</GID>
<name>OUT_1</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>208,-180.5,209,-180.5</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>208 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-168,199,-158</points>
<intersection>-168 4</intersection>
<intersection>-158 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>199,-158,203.5,-158</points>
<intersection>199 0</intersection>
<intersection>203.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>199,-168,215,-168</points>
<intersection>199 0</intersection>
<intersection>202.5 15</intersection>
<intersection>215 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>215,-168,215,-167.5</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<connection>
<GID>61</GID>
<name>clear</name></connection>
<intersection>-168 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>203.5,-158.5,203.5,-158</points>
<connection>
<GID>64</GID>
<name>count_enable</name></connection>
<intersection>-158 3</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>202.5,-168,202.5,-167.5</points>
<connection>
<GID>64</GID>
<name>clock</name></connection>
<intersection>-168 4</intersection></vsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240.5,-205,240.5,-188</points>
<connection>
<GID>74</GID>
<name>IN_3</name></connection>
<intersection>-201 1</intersection>
<intersection>-188 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235,-201,240.5,-201</points>
<intersection>235 17</intersection>
<intersection>240.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>239,-188,240.5,-188</points>
<connection>
<GID>75</GID>
<name>OUT_3</name></connection>
<intersection>240.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>235,-201,235,-200.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>-201 1</intersection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257,-168,257,-167.5</points>
<connection>
<GID>49</GID>
<name>clear</name></connection>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>-168 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>241,-168,257,-168</points>
<intersection>241 4</intersection>
<intersection>244.5 8</intersection>
<intersection>257 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>241,-168,241,-158</points>
<intersection>-168 3</intersection>
<intersection>-158 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>241,-158,245.5,-158</points>
<intersection>241 4</intersection>
<intersection>245.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>245.5,-158.5,245.5,-158</points>
<connection>
<GID>52</GID>
<name>count_enable</name></connection>
<intersection>-158 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>244.5,-168,244.5,-167.5</points>
<connection>
<GID>52</GID>
<name>clock</name></connection>
<intersection>-168 3</intersection></vsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246.5,-168,246.5,-167.5</points>
<connection>
<GID>52</GID>
<name>clear</name></connection>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<intersection>-167.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230.5,-167.5,246.5,-167.5</points>
<connection>
<GID>55</GID>
<name>clock</name></connection>
<intersection>230.5 4</intersection>
<intersection>246.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>230.5,-167.5,230.5,-158</points>
<intersection>-167.5 1</intersection>
<intersection>-158 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>230.5,-158,235,-158</points>
<intersection>230.5 4</intersection>
<intersection>235 17</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>235,-158.5,235,-158</points>
<connection>
<GID>55</GID>
<name>count_enable</name></connection>
<intersection>-158 15</intersection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,-208,239,-191</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>-208 5</intersection>
<intersection>-200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>237,-200.5,239,-200.5</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>239 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>239,-208,240.5,-208</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>239 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-206,240,-189</points>
<intersection>-206 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240,-206,240.5,-206</points>
<connection>
<GID>74</GID>
<name>IN_2</name></connection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>239,-189,240,-189</points>
<connection>
<GID>75</GID>
<name>OUT_2</name></connection>
<intersection>240 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239.5,-207,239.5,-190</points>
<intersection>-207 3</intersection>
<intersection>-190 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>239,-190,239.5,-190</points>
<connection>
<GID>75</GID>
<name>OUT_1</name></connection>
<intersection>239.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>239.5,-207,240.5,-207</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>239.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,-194.5,236,-194</points>
<connection>
<GID>75</GID>
<name>clear</name></connection>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<intersection>-194.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>220,-194.5,236,-194.5</points>
<intersection>220 2</intersection>
<intersection>223.5 10</intersection>
<intersection>236 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-194.5,220,-184.5</points>
<intersection>-194.5 1</intersection>
<intersection>-184.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>220,-184.5,224.5,-184.5</points>
<intersection>220 2</intersection>
<intersection>224.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>224.5,-185,224.5,-184.5</points>
<connection>
<GID>78</GID>
<name>count_enable</name></connection>
<intersection>-184.5 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>223.5,-194.5,223.5,-194</points>
<connection>
<GID>78</GID>
<name>clock</name></connection>
<intersection>-194.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,-205,230,-188</points>
<connection>
<GID>77</GID>
<name>IN_3</name></connection>
<intersection>-201 1</intersection>
<intersection>-188 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>224.5,-201,230,-201</points>
<intersection>224.5 17</intersection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228.5,-188,230,-188</points>
<connection>
<GID>78</GID>
<name>OUT_3</name></connection>
<intersection>230 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>224.5,-201,224.5,-200.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>-201 1</intersection></vsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,-208,228.5,-191</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>-208 5</intersection>
<intersection>-200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-200.5,228.5,-200.5</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>228.5,-208,230,-208</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>228.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,-206,229.5,-189</points>
<intersection>-206 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229.5,-206,230,-206</points>
<connection>
<GID>77</GID>
<name>IN_2</name></connection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228.5,-189,229.5,-189</points>
<connection>
<GID>78</GID>
<name>OUT_2</name></connection>
<intersection>229.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-207,229,-190</points>
<intersection>-207 3</intersection>
<intersection>-190 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>228.5,-190,229,-190</points>
<connection>
<GID>78</GID>
<name>OUT_1</name></connection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>229,-207,230,-207</points>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>229 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,-205,219.5,-188</points>
<connection>
<GID>80</GID>
<name>IN_3</name></connection>
<intersection>-201 1</intersection>
<intersection>-188 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>214,-201,219.5,-201</points>
<intersection>214 17</intersection>
<intersection>219.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>218,-188,219.5,-188</points>
<connection>
<GID>81</GID>
<name>OUT_3</name></connection>
<intersection>219.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>214,-201,214,-200.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>-201 1</intersection></vsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-208,218,-191</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<intersection>-208 5</intersection>
<intersection>-200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-200.5,218,-200.5</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>218,-208,219.5,-208</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-206,219,-189</points>
<intersection>-206 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,-206,219.5,-206</points>
<connection>
<GID>80</GID>
<name>IN_2</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>218,-189,219,-189</points>
<connection>
<GID>81</GID>
<name>OUT_2</name></connection>
<intersection>219 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-207,218.5,-190</points>
<intersection>-207 3</intersection>
<intersection>-190 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>218,-190,218.5,-190</points>
<connection>
<GID>81</GID>
<name>OUT_1</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>218.5,-207,219.5,-207</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>218.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209.5,-194,209.5,-184.5</points>
<intersection>-194 4</intersection>
<intersection>-184.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>209.5,-184.5,214,-184.5</points>
<intersection>209.5 0</intersection>
<intersection>214 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>209.5,-194,225.5,-194</points>
<connection>
<GID>81</GID>
<name>clock</name></connection>
<intersection>209.5 0</intersection>
<intersection>225.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>225.5,-194.5,225.5,-194</points>
<connection>
<GID>78</GID>
<name>clear</name></connection>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>-194 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>214,-185,214,-184.5</points>
<connection>
<GID>81</GID>
<name>count_enable</name></connection>
<intersection>-184.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209,-205,209,-188</points>
<connection>
<GID>83</GID>
<name>IN_3</name></connection>
<intersection>-201 1</intersection>
<intersection>-188 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203.5,-201,209,-201</points>
<intersection>203.5 17</intersection>
<intersection>209 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207.5,-188,209,-188</points>
<connection>
<GID>84</GID>
<name>OUT_3</name></connection>
<intersection>209 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>203.5,-201,203.5,-200.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>-201 1</intersection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,-208,207.5,-191</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>-208 5</intersection>
<intersection>-200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>205.5,-200.5,207.5,-200.5</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>207.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>207.5,-208,209,-208</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>207.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-206,208.5,-189</points>
<intersection>-206 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208.5,-206,209,-206</points>
<connection>
<GID>83</GID>
<name>IN_2</name></connection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207.5,-189,208.5,-189</points>
<connection>
<GID>84</GID>
<name>OUT_2</name></connection>
<intersection>208.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-207,208,-190</points>
<intersection>-207 3</intersection>
<intersection>-190 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>207.5,-190,208,-190</points>
<connection>
<GID>84</GID>
<name>OUT_1</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>208,-207,209,-207</points>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<intersection>208 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-194.5,199,-184.5</points>
<intersection>-194.5 4</intersection>
<intersection>-184.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>199,-184.5,203.5,-184.5</points>
<intersection>199 0</intersection>
<intersection>203.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>199,-194.5,215,-194.5</points>
<intersection>199 0</intersection>
<intersection>202.5 15</intersection>
<intersection>215 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>215,-194.5,215,-194</points>
<connection>
<GID>81</GID>
<name>clear</name></connection>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<intersection>-194.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>203.5,-185,203.5,-184.5</points>
<connection>
<GID>84</GID>
<name>count_enable</name></connection>
<intersection>-184.5 3</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>202.5,-194.5,202.5,-194</points>
<connection>
<GID>84</GID>
<name>clock</name></connection>
<intersection>-194.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257,-194.5,257,-194</points>
<connection>
<GID>69</GID>
<name>clear</name></connection>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>-194.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>241,-194.5,257,-194.5</points>
<intersection>241 4</intersection>
<intersection>244.5 8</intersection>
<intersection>257 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>241,-194.5,241,-184.5</points>
<intersection>-194.5 3</intersection>
<intersection>-184.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>241,-184.5,245.5,-184.5</points>
<intersection>241 4</intersection>
<intersection>245.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>245.5,-185,245.5,-184.5</points>
<connection>
<GID>72</GID>
<name>count_enable</name></connection>
<intersection>-184.5 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>244.5,-194.5,244.5,-194</points>
<connection>
<GID>72</GID>
<name>clock</name></connection>
<intersection>-194.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246.5,-194.5,246.5,-194</points>
<connection>
<GID>72</GID>
<name>clear</name></connection>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<intersection>-194.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230.5,-194.5,246.5,-194.5</points>
<intersection>230.5 4</intersection>
<intersection>234 20</intersection>
<intersection>246.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>230.5,-194.5,230.5,-185</points>
<intersection>-194.5 1</intersection>
<intersection>-185 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>230.5,-185,235,-185</points>
<connection>
<GID>75</GID>
<name>count_enable</name></connection>
<intersection>230.5 4</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>234,-194.5,234,-194</points>
<connection>
<GID>75</GID>
<name>clock</name></connection>
<intersection>-194.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303,-151,303,-134</points>
<connection>
<GID>86</GID>
<name>IN_3</name></connection>
<intersection>-147 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>297.5,-147,303,-147</points>
<intersection>297.5 17</intersection>
<intersection>303 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301.5,-134,303,-134</points>
<connection>
<GID>87</GID>
<name>OUT_3</name></connection>
<intersection>303 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>297.5,-147,297.5,-146.5</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>-147 1</intersection></vsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-154,301.5,-137</points>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection>
<intersection>-154 5</intersection>
<intersection>-146.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>299.5,-146.5,301.5,-146.5</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>301.5,-154,303,-154</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,-152,302.5,-135</points>
<intersection>-152 1</intersection>
<intersection>-135 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302.5,-152,303,-152</points>
<connection>
<GID>86</GID>
<name>IN_2</name></connection>
<intersection>302.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301.5,-135,302.5,-135</points>
<connection>
<GID>87</GID>
<name>OUT_2</name></connection>
<intersection>302.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-153,302,-136</points>
<intersection>-153 3</intersection>
<intersection>-136 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>301.5,-136,302,-136</points>
<connection>
<GID>87</GID>
<name>OUT_1</name></connection>
<intersection>302 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>302,-153,303,-153</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>302 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298.5,-140.5,298.5,-140</points>
<connection>
<GID>88</GID>
<name>OUT</name></connection>
<connection>
<GID>87</GID>
<name>clear</name></connection>
<intersection>-140.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282.5,-140.5,298.5,-140.5</points>
<intersection>282.5 2</intersection>
<intersection>286 7</intersection>
<intersection>298.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>282.5,-140.5,282.5,-130.5</points>
<intersection>-140.5 1</intersection>
<intersection>-130.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>282.5,-130.5,287,-130.5</points>
<intersection>282.5 2</intersection>
<intersection>287 10</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>286,-140.5,286,-140</points>
<connection>
<GID>90</GID>
<name>clock</name></connection>
<intersection>-140.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>287,-131,287,-130.5</points>
<connection>
<GID>90</GID>
<name>count_enable</name></connection>
<intersection>-130.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,-151,292.5,-134</points>
<connection>
<GID>89</GID>
<name>IN_3</name></connection>
<intersection>-147 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287,-147,292.5,-147</points>
<intersection>287 17</intersection>
<intersection>292.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>291,-134,292.5,-134</points>
<connection>
<GID>90</GID>
<name>OUT_3</name></connection>
<intersection>292.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>287,-147,287,-146.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>-147 1</intersection></vsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,-154,291,-137</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<intersection>-154 5</intersection>
<intersection>-146.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>289,-146.5,291,-146.5</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>291 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>291,-154,292.5,-154</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>291 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,-152,292,-135</points>
<intersection>-152 1</intersection>
<intersection>-135 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>292,-152,292.5,-152</points>
<connection>
<GID>89</GID>
<name>IN_2</name></connection>
<intersection>292 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>291,-135,292,-135</points>
<connection>
<GID>90</GID>
<name>OUT_2</name></connection>
<intersection>292 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,-153,291.5,-136</points>
<intersection>-153 3</intersection>
<intersection>-136 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>291,-136,291.5,-136</points>
<connection>
<GID>90</GID>
<name>OUT_1</name></connection>
<intersection>291.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>291.5,-153,292.5,-153</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,-140.5,288,-140</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<connection>
<GID>90</GID>
<name>clear</name></connection>
<intersection>-140.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>272,-140.5,288,-140.5</points>
<intersection>272 2</intersection>
<intersection>275.5 12</intersection>
<intersection>288 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>272,-140.5,272,-131</points>
<intersection>-140.5 1</intersection>
<intersection>-131 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>272,-131,276.5,-131</points>
<connection>
<GID>93</GID>
<name>count_enable</name></connection>
<intersection>272 2</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>275.5,-140.5,275.5,-140</points>
<connection>
<GID>93</GID>
<name>clock</name></connection>
<intersection>-140.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-151,282,-134</points>
<connection>
<GID>92</GID>
<name>IN_3</name></connection>
<intersection>-147 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276.5,-147,282,-147</points>
<intersection>276.5 17</intersection>
<intersection>282 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280.5,-134,282,-134</points>
<connection>
<GID>93</GID>
<name>OUT_3</name></connection>
<intersection>282 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>276.5,-147,276.5,-146.5</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>-147 1</intersection></vsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280.5,-154,280.5,-137</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<intersection>-154 5</intersection>
<intersection>-146.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>278.5,-146.5,280.5,-146.5</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>280.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>280.5,-154,282,-154</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>280.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-152,281.5,-135</points>
<intersection>-152 1</intersection>
<intersection>-135 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281.5,-152,282,-152</points>
<connection>
<GID>92</GID>
<name>IN_2</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280.5,-135,281.5,-135</points>
<connection>
<GID>93</GID>
<name>OUT_2</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,-153,281,-136</points>
<intersection>-153 3</intersection>
<intersection>-136 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>280.5,-136,281,-136</points>
<connection>
<GID>93</GID>
<name>OUT_1</name></connection>
<intersection>281 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>281,-153,282,-153</points>
<connection>
<GID>92</GID>
<name>IN_1</name></connection>
<intersection>281 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,-151,271.5,-134</points>
<connection>
<GID>95</GID>
<name>IN_3</name></connection>
<intersection>-147 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266,-147,271.5,-147</points>
<intersection>266 17</intersection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>270,-134,271.5,-134</points>
<connection>
<GID>126</GID>
<name>OUT_3</name></connection>
<intersection>271.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>266,-147,266,-146.5</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>-147 1</intersection></vsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,-154,270,-137</points>
<connection>
<GID>126</GID>
<name>OUT_0</name></connection>
<intersection>-154 5</intersection>
<intersection>-146.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>268,-146.5,270,-146.5</points>
<connection>
<GID>127</GID>
<name>IN_1</name></connection>
<intersection>270 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>270,-154,271.5,-154</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>270 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-152,271,-135</points>
<intersection>-152 1</intersection>
<intersection>-135 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>271,-152,271.5,-152</points>
<connection>
<GID>95</GID>
<name>IN_2</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>270,-135,271,-135</points>
<connection>
<GID>126</GID>
<name>OUT_2</name></connection>
<intersection>271 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-153,270.5,-136</points>
<intersection>-153 3</intersection>
<intersection>-136 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>270,-136,270.5,-136</points>
<connection>
<GID>126</GID>
<name>OUT_1</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>270.5,-153,271.5,-153</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,-140.5,261.5,-130.5</points>
<intersection>-140.5 4</intersection>
<intersection>-130.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>261.5,-130.5,266,-130.5</points>
<intersection>261.5 0</intersection>
<intersection>266 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>261.5,-140.5,277.5,-140.5</points>
<intersection>261.5 0</intersection>
<intersection>265 7</intersection>
<intersection>277.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>277.5,-140.5,277.5,-140</points>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<connection>
<GID>93</GID>
<name>clear</name></connection>
<intersection>-140.5 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>265,-140.5,265,-140</points>
<connection>
<GID>126</GID>
<name>clock</name></connection>
<intersection>-140.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>266,-131,266,-130.5</points>
<connection>
<GID>126</GID>
<name>count_enable</name></connection>
<intersection>-130.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,-151,261,-134</points>
<connection>
<GID>128</GID>
<name>IN_3</name></connection>
<intersection>-147 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255.5,-147,261,-147</points>
<intersection>255.5 17</intersection>
<intersection>261 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259.5,-134,261,-134</points>
<connection>
<GID>129</GID>
<name>OUT_3</name></connection>
<intersection>261 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>255.5,-147,255.5,-146.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>-147 1</intersection></vsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,-154,259.5,-137</points>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<intersection>-154 5</intersection>
<intersection>-146.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>257.5,-146.5,259.5,-146.5</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>259.5,-154,261,-154</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>259.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,-152,260.5,-135</points>
<intersection>-152 1</intersection>
<intersection>-135 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,-152,261,-152</points>
<connection>
<GID>128</GID>
<name>IN_2</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259.5,-135,260.5,-135</points>
<connection>
<GID>129</GID>
<name>OUT_2</name></connection>
<intersection>260.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-153,260,-136</points>
<intersection>-153 3</intersection>
<intersection>-136 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>259.5,-136,260,-136</points>
<connection>
<GID>129</GID>
<name>OUT_1</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>260,-153,261,-153</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,-140,251,-130.5</points>
<intersection>-140 4</intersection>
<intersection>-130.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>251,-130.5,255.5,-130.5</points>
<intersection>251 0</intersection>
<intersection>255.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>251,-140,267,-140</points>
<connection>
<GID>129</GID>
<name>clock</name></connection>
<intersection>251 0</intersection>
<intersection>267 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>267,-140.5,267,-140</points>
<connection>
<GID>127</GID>
<name>OUT</name></connection>
<connection>
<GID>126</GID>
<name>clear</name></connection>
<intersection>-140 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>255.5,-131,255.5,-130.5</points>
<connection>
<GID>129</GID>
<name>count_enable</name></connection>
<intersection>-130.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-140,293,-130</points>
<intersection>-140 4</intersection>
<intersection>-130 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>197.5,-130,297.5,-130</points>
<intersection>197.5 7</intersection>
<intersection>293 0</intersection>
<intersection>297.5 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293,-140,296.5,-140</points>
<connection>
<GID>87</GID>
<name>clock</name></connection>
<intersection>293 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>297.5,-131,297.5,-130</points>
<connection>
<GID>87</GID>
<name>count_enable</name></connection>
<intersection>-130 3</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>197.5,-167.5,197.5,-130</points>
<intersection>-167.5 8</intersection>
<intersection>-130 3</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>197.5,-167.5,204.5,-167.5</points>
<connection>
<GID>64</GID>
<name>clear</name></connection>
<intersection>197.5 7</intersection>
<intersection>204.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>204.5,-168,204.5,-167.5</points>
<connection>
<GID>65</GID>
<name>OUT</name></connection>
<intersection>-167.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,-151,250.5,-134</points>
<connection>
<GID>131</GID>
<name>IN_3</name></connection>
<intersection>-147 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245,-147,250.5,-147</points>
<intersection>245 17</intersection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>249,-134,250.5,-134</points>
<connection>
<GID>132</GID>
<name>OUT_3</name></connection>
<intersection>250.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>245,-147,245,-146.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>-147 1</intersection></vsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303,-124.5,303,-107.5</points>
<connection>
<GID>96</GID>
<name>IN_3</name></connection>
<intersection>-120.5 1</intersection>
<intersection>-107.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>297.5,-120.5,303,-120.5</points>
<intersection>297.5 17</intersection>
<intersection>303 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301.5,-107.5,303,-107.5</points>
<connection>
<GID>97</GID>
<name>OUT_3</name></connection>
<intersection>303 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>297.5,-120.5,297.5,-120</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>-120.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-127.5,301.5,-110.5</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>-127.5 5</intersection>
<intersection>-120 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>299.5,-120,301.5,-120</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>301.5,-127.5,303,-127.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,-125.5,302.5,-108.5</points>
<intersection>-125.5 1</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302.5,-125.5,303,-125.5</points>
<connection>
<GID>96</GID>
<name>IN_2</name></connection>
<intersection>302.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301.5,-108.5,302.5,-108.5</points>
<connection>
<GID>97</GID>
<name>OUT_2</name></connection>
<intersection>302.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-126.5,302,-109.5</points>
<intersection>-126.5 3</intersection>
<intersection>-109.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>301.5,-109.5,302,-109.5</points>
<connection>
<GID>97</GID>
<name>OUT_1</name></connection>
<intersection>302 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>302,-126.5,303,-126.5</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>302 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298.5,-114,298.5,-113.5</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<connection>
<GID>97</GID>
<name>clear</name></connection>
<intersection>-114 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282.5,-114,298.5,-114</points>
<intersection>282.5 2</intersection>
<intersection>286 7</intersection>
<intersection>298.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>282.5,-114,282.5,-104</points>
<intersection>-114 1</intersection>
<intersection>-104 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>282.5,-104,287,-104</points>
<intersection>282.5 2</intersection>
<intersection>287 10</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>286,-114,286,-113.5</points>
<connection>
<GID>100</GID>
<name>clock</name></connection>
<intersection>-114 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>287,-104.5,287,-104</points>
<connection>
<GID>100</GID>
<name>count_enable</name></connection>
<intersection>-104 5</intersection></vsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249,-154,249,-137</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>-154 5</intersection>
<intersection>-146.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>247,-146.5,249,-146.5</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<intersection>249 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>249,-154,250.5,-154</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>249 0</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,-124.5,292.5,-107.5</points>
<connection>
<GID>99</GID>
<name>IN_3</name></connection>
<intersection>-120.5 1</intersection>
<intersection>-107.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287,-120.5,292.5,-120.5</points>
<intersection>287 17</intersection>
<intersection>292.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>291,-107.5,292.5,-107.5</points>
<connection>
<GID>100</GID>
<name>OUT_3</name></connection>
<intersection>292.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>287,-120.5,287,-120</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-120.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,-127.5,291,-110.5</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<intersection>-127.5 5</intersection>
<intersection>-120 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>289,-120,291,-120</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>291 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>291,-127.5,292.5,-127.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>291 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,-125.5,292,-108.5</points>
<intersection>-125.5 1</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>292,-125.5,292.5,-125.5</points>
<connection>
<GID>99</GID>
<name>IN_2</name></connection>
<intersection>292 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>291,-108.5,292,-108.5</points>
<connection>
<GID>100</GID>
<name>OUT_2</name></connection>
<intersection>292 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,-126.5,291.5,-109.5</points>
<intersection>-126.5 3</intersection>
<intersection>-109.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>291,-109.5,291.5,-109.5</points>
<connection>
<GID>100</GID>
<name>OUT_1</name></connection>
<intersection>291.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>291.5,-126.5,292.5,-126.5</points>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,-114,288,-113.5</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<connection>
<GID>100</GID>
<name>clear</name></connection>
<intersection>-113.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>272,-113.5,288,-113.5</points>
<connection>
<GID>103</GID>
<name>clock</name></connection>
<intersection>272 2</intersection>
<intersection>288 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>272,-113.5,272,-104</points>
<intersection>-113.5 1</intersection>
<intersection>-104 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>272,-104,276.5,-104</points>
<intersection>272 2</intersection>
<intersection>276.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>276.5,-104.5,276.5,-104</points>
<connection>
<GID>103</GID>
<name>count_enable</name></connection>
<intersection>-104 5</intersection></vsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-124.5,282,-107.5</points>
<connection>
<GID>102</GID>
<name>IN_3</name></connection>
<intersection>-120.5 1</intersection>
<intersection>-107.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276.5,-120.5,282,-120.5</points>
<intersection>276.5 17</intersection>
<intersection>282 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280.5,-107.5,282,-107.5</points>
<connection>
<GID>103</GID>
<name>OUT_3</name></connection>
<intersection>282 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>276.5,-120.5,276.5,-120</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>-120.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280.5,-127.5,280.5,-110.5</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<intersection>-127.5 5</intersection>
<intersection>-120 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>278.5,-120,280.5,-120</points>
<connection>
<GID>104</GID>
<name>IN_1</name></connection>
<intersection>280.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>280.5,-127.5,282,-127.5</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>280.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-125.5,281.5,-108.5</points>
<intersection>-125.5 1</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281.5,-125.5,282,-125.5</points>
<connection>
<GID>102</GID>
<name>IN_2</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280.5,-108.5,281.5,-108.5</points>
<connection>
<GID>103</GID>
<name>OUT_2</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,-126.5,281,-109.5</points>
<intersection>-126.5 3</intersection>
<intersection>-109.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>280.5,-109.5,281,-109.5</points>
<connection>
<GID>103</GID>
<name>OUT_1</name></connection>
<intersection>281 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>281,-126.5,282,-126.5</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>281 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,-124.5,271.5,-107.5</points>
<connection>
<GID>105</GID>
<name>IN_3</name></connection>
<intersection>-120.5 1</intersection>
<intersection>-107.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266,-120.5,271.5,-120.5</points>
<intersection>266 17</intersection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>270,-107.5,271.5,-107.5</points>
<connection>
<GID>106</GID>
<name>OUT_3</name></connection>
<intersection>271.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>266,-120.5,266,-120</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>-120.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,-127.5,270,-110.5</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>-127.5 5</intersection>
<intersection>-120 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>268,-120,270,-120</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>270 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>270,-127.5,271.5,-127.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>270 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-125.5,271,-108.5</points>
<intersection>-125.5 1</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>271,-125.5,271.5,-125.5</points>
<connection>
<GID>105</GID>
<name>IN_2</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>270,-108.5,271,-108.5</points>
<connection>
<GID>106</GID>
<name>OUT_2</name></connection>
<intersection>271 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-126.5,270.5,-109.5</points>
<intersection>-126.5 3</intersection>
<intersection>-109.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>270,-109.5,270.5,-109.5</points>
<connection>
<GID>106</GID>
<name>OUT_1</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>270.5,-126.5,271.5,-126.5</points>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,-114,261.5,-104</points>
<intersection>-114 4</intersection>
<intersection>-104 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>261.5,-104,266,-104</points>
<intersection>261.5 0</intersection>
<intersection>266 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>261.5,-114,277.5,-114</points>
<intersection>261.5 0</intersection>
<intersection>265 7</intersection>
<intersection>277.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>277.5,-114,277.5,-113.5</points>
<connection>
<GID>104</GID>
<name>OUT</name></connection>
<connection>
<GID>103</GID>
<name>clear</name></connection>
<intersection>-114 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>265,-114,265,-113.5</points>
<connection>
<GID>106</GID>
<name>clock</name></connection>
<intersection>-114 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>266,-104.5,266,-104</points>
<connection>
<GID>106</GID>
<name>count_enable</name></connection>
<intersection>-104 3</intersection></vsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,-124.5,261,-107.5</points>
<connection>
<GID>108</GID>
<name>IN_3</name></connection>
<intersection>-120.5 1</intersection>
<intersection>-107.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255.5,-120.5,261,-120.5</points>
<intersection>255.5 17</intersection>
<intersection>261 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259.5,-107.5,261,-107.5</points>
<connection>
<GID>109</GID>
<name>OUT_3</name></connection>
<intersection>261 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>255.5,-120.5,255.5,-120</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>-120.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,-127.5,259.5,-110.5</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<intersection>-127.5 5</intersection>
<intersection>-120 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>257.5,-120,259.5,-120</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>259.5,-127.5,261,-127.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>259.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,-125.5,260.5,-108.5</points>
<intersection>-125.5 1</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,-125.5,261,-125.5</points>
<connection>
<GID>108</GID>
<name>IN_2</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259.5,-108.5,260.5,-108.5</points>
<connection>
<GID>109</GID>
<name>OUT_2</name></connection>
<intersection>260.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-126.5,260,-109.5</points>
<intersection>-126.5 3</intersection>
<intersection>-109.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>259.5,-109.5,260,-109.5</points>
<connection>
<GID>109</GID>
<name>OUT_1</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>260,-126.5,261,-126.5</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,-152,250,-135</points>
<intersection>-152 1</intersection>
<intersection>-135 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250,-152,250.5,-152</points>
<connection>
<GID>131</GID>
<name>IN_2</name></connection>
<intersection>250 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>249,-135,250,-135</points>
<connection>
<GID>132</GID>
<name>OUT_2</name></connection>
<intersection>250 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,-113.5,251,-104</points>
<intersection>-113.5 4</intersection>
<intersection>-104 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>251,-104,255.5,-104</points>
<intersection>251 0</intersection>
<intersection>255.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>251,-113.5,267,-113.5</points>
<connection>
<GID>109</GID>
<name>clock</name></connection>
<intersection>251 0</intersection>
<intersection>267 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>267,-114,267,-113.5</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<connection>
<GID>106</GID>
<name>clear</name></connection>
<intersection>-113.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>255.5,-104.5,255.5,-104</points>
<connection>
<GID>109</GID>
<name>count_enable</name></connection>
<intersection>-104 3</intersection></vsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-113.5,293,-104</points>
<intersection>-113.5 4</intersection>
<intersection>-104 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>293,-104,297.5,-104</points>
<intersection>293 0</intersection>
<intersection>297.5 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293,-113.5,296.5,-113.5</points>
<connection>
<GID>97</GID>
<name>clock</name></connection>
<intersection>293 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>297.5,-104.5,297.5,-103</points>
<connection>
<GID>97</GID>
<name>count_enable</name></connection>
<intersection>-104 3</intersection>
<intersection>-103 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>196.5,-103,297.5,-103</points>
<intersection>196.5 7</intersection>
<intersection>297.5 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>196.5,-140.5,196.5,-103</points>
<intersection>-140.5 8</intersection>
<intersection>-103 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>196.5,-140.5,204,-140.5</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<intersection>196.5 7</intersection>
<intersection>204 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>204,-140.5,204,-140</points>
<connection>
<GID>144</GID>
<name>clear</name></connection>
<intersection>-140.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,-124.5,250.5,-107.5</points>
<connection>
<GID>111</GID>
<name>IN_3</name></connection>
<intersection>-120.5 1</intersection>
<intersection>-107.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245,-120.5,250.5,-120.5</points>
<intersection>245 17</intersection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>249,-107.5,250.5,-107.5</points>
<connection>
<GID>112</GID>
<name>OUT_3</name></connection>
<intersection>250.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>245,-120.5,245,-120</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>-120.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249,-127.5,249,-110.5</points>
<connection>
<GID>112</GID>
<name>OUT_0</name></connection>
<intersection>-127.5 5</intersection>
<intersection>-120 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>247,-120,249,-120</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>249 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>249,-127.5,250.5,-127.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>249 0</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,-125.5,250,-108.5</points>
<intersection>-125.5 1</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250,-125.5,250.5,-125.5</points>
<connection>
<GID>111</GID>
<name>IN_2</name></connection>
<intersection>250 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>249,-108.5,250,-108.5</points>
<connection>
<GID>112</GID>
<name>OUT_2</name></connection>
<intersection>250 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,-126.5,249.5,-109.5</points>
<intersection>-126.5 3</intersection>
<intersection>-109.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>249,-109.5,249.5,-109.5</points>
<connection>
<GID>112</GID>
<name>OUT_1</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>249.5,-126.5,250.5,-126.5</points>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<intersection>249.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,-153,249.5,-136</points>
<intersection>-153 3</intersection>
<intersection>-136 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>249,-136,249.5,-136</points>
<connection>
<GID>132</GID>
<name>OUT_1</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>249.5,-153,250.5,-153</points>
<connection>
<GID>131</GID>
<name>IN_1</name></connection>
<intersection>249.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-124.5,240,-107.5</points>
<connection>
<GID>114</GID>
<name>IN_3</name></connection>
<intersection>-120.5 1</intersection>
<intersection>-107.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234.5,-120.5,240,-120.5</points>
<intersection>234.5 17</intersection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-107.5,240,-107.5</points>
<connection>
<GID>115</GID>
<name>OUT_3</name></connection>
<intersection>240 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>234.5,-120.5,234.5,-120</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>-120.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,-127.5,238.5,-110.5</points>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<intersection>-127.5 5</intersection>
<intersection>-120 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>236.5,-120,238.5,-120</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>238.5,-127.5,240,-127.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>238.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239.5,-125.5,239.5,-108.5</points>
<intersection>-125.5 1</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239.5,-125.5,240,-125.5</points>
<connection>
<GID>114</GID>
<name>IN_2</name></connection>
<intersection>239.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-108.5,239.5,-108.5</points>
<connection>
<GID>115</GID>
<name>OUT_2</name></connection>
<intersection>239.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,-126.5,239,-109.5</points>
<intersection>-126.5 3</intersection>
<intersection>-109.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-109.5,239,-109.5</points>
<connection>
<GID>115</GID>
<name>OUT_1</name></connection>
<intersection>239 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>239,-126.5,240,-126.5</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>239 0</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235.5,-114,235.5,-113.5</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<connection>
<GID>115</GID>
<name>clear</name></connection>
<intersection>-114 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219.5,-114,235.5,-114</points>
<intersection>219.5 2</intersection>
<intersection>223 10</intersection>
<intersection>235.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>219.5,-114,219.5,-104</points>
<intersection>-114 1</intersection>
<intersection>-104 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>219.5,-104,224,-104</points>
<intersection>219.5 2</intersection>
<intersection>224 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>224,-104.5,224,-104</points>
<connection>
<GID>118</GID>
<name>count_enable</name></connection>
<intersection>-104 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>223,-114,223,-113.5</points>
<connection>
<GID>118</GID>
<name>clock</name></connection>
<intersection>-114 1</intersection></vsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,-124.5,229.5,-107.5</points>
<connection>
<GID>117</GID>
<name>IN_3</name></connection>
<intersection>-120.5 1</intersection>
<intersection>-107.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>224,-120.5,229.5,-120.5</points>
<intersection>224 17</intersection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228,-107.5,229.5,-107.5</points>
<connection>
<GID>118</GID>
<name>OUT_3</name></connection>
<intersection>229.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>224,-120.5,224,-120</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-120.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,-127.5,228,-110.5</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<intersection>-127.5 5</intersection>
<intersection>-120 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-120,228,-120</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>228 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>228,-127.5,229.5,-127.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>228 0</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-125.5,229,-108.5</points>
<intersection>-125.5 1</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229,-125.5,229.5,-125.5</points>
<connection>
<GID>117</GID>
<name>IN_2</name></connection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228,-108.5,229,-108.5</points>
<connection>
<GID>118</GID>
<name>OUT_2</name></connection>
<intersection>229 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,-126.5,228.5,-109.5</points>
<intersection>-126.5 3</intersection>
<intersection>-109.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>228,-109.5,228.5,-109.5</points>
<connection>
<GID>118</GID>
<name>OUT_1</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>228.5,-126.5,229.5,-126.5</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>228.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-124.5,219,-107.5</points>
<connection>
<GID>120</GID>
<name>IN_3</name></connection>
<intersection>-120.5 1</intersection>
<intersection>-107.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213.5,-120.5,219,-120.5</points>
<intersection>213.5 17</intersection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>217.5,-107.5,219,-107.5</points>
<connection>
<GID>121</GID>
<name>OUT_3</name></connection>
<intersection>219 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>213.5,-120.5,213.5,-120</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>-120.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217.5,-127.5,217.5,-110.5</points>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection>
<intersection>-127.5 5</intersection>
<intersection>-120 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>215.5,-120,217.5,-120</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>217.5,-127.5,219,-127.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-125.5,218.5,-108.5</points>
<intersection>-125.5 1</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218.5,-125.5,219,-125.5</points>
<connection>
<GID>120</GID>
<name>IN_2</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>217.5,-108.5,218.5,-108.5</points>
<connection>
<GID>121</GID>
<name>OUT_2</name></connection>
<intersection>218.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-126.5,218,-109.5</points>
<intersection>-126.5 3</intersection>
<intersection>-109.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>217.5,-109.5,218,-109.5</points>
<connection>
<GID>121</GID>
<name>OUT_1</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>218,-126.5,219,-126.5</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209,-113.5,209,-104</points>
<intersection>-113.5 4</intersection>
<intersection>-104 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>209,-104,213.5,-104</points>
<intersection>209 0</intersection>
<intersection>213.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>209,-113.5,225,-113.5</points>
<connection>
<GID>121</GID>
<name>clock</name></connection>
<intersection>209 0</intersection>
<intersection>225 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>225,-114,225,-113.5</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<connection>
<GID>118</GID>
<name>clear</name></connection>
<intersection>-113.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>213.5,-104.5,213.5,-104</points>
<connection>
<GID>121</GID>
<name>count_enable</name></connection>
<intersection>-104 3</intersection></vsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-124.5,208.5,-107.5</points>
<connection>
<GID>123</GID>
<name>IN_3</name></connection>
<intersection>-120.5 1</intersection>
<intersection>-107.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-120.5,208.5,-120.5</points>
<intersection>203 17</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207,-107.5,208.5,-107.5</points>
<connection>
<GID>124</GID>
<name>OUT_3</name></connection>
<intersection>208.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>203,-120.5,203,-120</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>-120.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-127.5,207,-110.5</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>-127.5 5</intersection>
<intersection>-120 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>205,-120,207,-120</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>207,-127.5,208.5,-127.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-125.5,208,-108.5</points>
<intersection>-125.5 1</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208,-125.5,208.5,-125.5</points>
<connection>
<GID>123</GID>
<name>IN_2</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207,-108.5,208,-108.5</points>
<connection>
<GID>124</GID>
<name>OUT_2</name></connection>
<intersection>208 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,-126.5,207.5,-109.5</points>
<intersection>-126.5 3</intersection>
<intersection>-109.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>207,-109.5,207.5,-109.5</points>
<connection>
<GID>124</GID>
<name>OUT_1</name></connection>
<intersection>207.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>207.5,-126.5,208.5,-126.5</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<intersection>207.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-114,198.5,-104</points>
<intersection>-114 4</intersection>
<intersection>-104 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198.5,-104,203,-104</points>
<intersection>198.5 0</intersection>
<intersection>203 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>198.5,-114,214.5,-114</points>
<intersection>198.5 0</intersection>
<intersection>202 15</intersection>
<intersection>214.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>214.5,-114,214.5,-113.5</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<connection>
<GID>121</GID>
<name>clear</name></connection>
<intersection>-114 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>203,-104.5,203,-104</points>
<connection>
<GID>124</GID>
<name>count_enable</name></connection>
<intersection>-104 3</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>202,-114,202,-113.5</points>
<connection>
<GID>124</GID>
<name>clock</name></connection>
<intersection>-114 4</intersection></vsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-151,240,-134</points>
<connection>
<GID>134</GID>
<name>IN_3</name></connection>
<intersection>-147 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234.5,-147,240,-147</points>
<intersection>234.5 17</intersection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-134,240,-134</points>
<connection>
<GID>135</GID>
<name>OUT_3</name></connection>
<intersection>240 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>234.5,-147,234.5,-146.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-147 1</intersection></vsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>256.5,-114,256.5,-113.5</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<connection>
<GID>109</GID>
<name>clear</name></connection>
<intersection>-114 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>240.5,-114,256.5,-114</points>
<intersection>240.5 4</intersection>
<intersection>244 8</intersection>
<intersection>256.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>240.5,-114,240.5,-104</points>
<intersection>-114 3</intersection>
<intersection>-104 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>240.5,-104,245,-104</points>
<intersection>240.5 4</intersection>
<intersection>245 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>245,-104.5,245,-104</points>
<connection>
<GID>112</GID>
<name>count_enable</name></connection>
<intersection>-104 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>244,-114,244,-113.5</points>
<connection>
<GID>112</GID>
<name>clock</name></connection>
<intersection>-114 3</intersection></vsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-114,246,-113.5</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<connection>
<GID>112</GID>
<name>clear</name></connection>
<intersection>-113.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230,-113.5,246,-113.5</points>
<connection>
<GID>115</GID>
<name>clock</name></connection>
<intersection>230 4</intersection>
<intersection>246 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>230,-113.5,230,-104</points>
<intersection>-113.5 1</intersection>
<intersection>-104 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>230,-104,234.5,-104</points>
<intersection>230 4</intersection>
<intersection>234.5 17</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>234.5,-104.5,234.5,-104</points>
<connection>
<GID>115</GID>
<name>count_enable</name></connection>
<intersection>-104 15</intersection></vsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,-154,238.5,-137</points>
<connection>
<GID>135</GID>
<name>OUT_0</name></connection>
<intersection>-154 5</intersection>
<intersection>-146.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>236.5,-146.5,238.5,-146.5</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>238.5,-154,240,-154</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>238.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239.5,-152,239.5,-135</points>
<intersection>-152 1</intersection>
<intersection>-135 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239.5,-152,240,-152</points>
<connection>
<GID>134</GID>
<name>IN_2</name></connection>
<intersection>239.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-135,239.5,-135</points>
<connection>
<GID>135</GID>
<name>OUT_2</name></connection>
<intersection>239.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,-153,239,-136</points>
<intersection>-153 3</intersection>
<intersection>-136 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-136,239,-136</points>
<connection>
<GID>135</GID>
<name>OUT_1</name></connection>
<intersection>239 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>239,-153,240,-153</points>
<connection>
<GID>134</GID>
<name>IN_1</name></connection>
<intersection>239 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235.5,-140.5,235.5,-140</points>
<connection>
<GID>136</GID>
<name>OUT</name></connection>
<connection>
<GID>135</GID>
<name>clear</name></connection>
<intersection>-140.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219.5,-140.5,235.5,-140.5</points>
<intersection>219.5 2</intersection>
<intersection>223 10</intersection>
<intersection>235.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>219.5,-140.5,219.5,-130.5</points>
<intersection>-140.5 1</intersection>
<intersection>-130.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>219.5,-130.5,224,-130.5</points>
<intersection>219.5 2</intersection>
<intersection>224 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>224,-131,224,-130.5</points>
<connection>
<GID>138</GID>
<name>count_enable</name></connection>
<intersection>-130.5 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>223,-140.5,223,-140</points>
<connection>
<GID>138</GID>
<name>clock</name></connection>
<intersection>-140.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,-151,229.5,-134</points>
<connection>
<GID>137</GID>
<name>IN_3</name></connection>
<intersection>-147 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>224,-147,229.5,-147</points>
<intersection>224 17</intersection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228,-134,229.5,-134</points>
<connection>
<GID>138</GID>
<name>OUT_3</name></connection>
<intersection>229.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>224,-147,224,-146.5</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>-147 1</intersection></vsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,-154,228,-137</points>
<connection>
<GID>138</GID>
<name>OUT_0</name></connection>
<intersection>-154 5</intersection>
<intersection>-146.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-146.5,228,-146.5</points>
<connection>
<GID>139</GID>
<name>IN_1</name></connection>
<intersection>228 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>228,-154,229.5,-154</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>228 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-152,229,-135</points>
<intersection>-152 1</intersection>
<intersection>-135 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229,-152,229.5,-152</points>
<connection>
<GID>137</GID>
<name>IN_2</name></connection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228,-135,229,-135</points>
<connection>
<GID>138</GID>
<name>OUT_2</name></connection>
<intersection>229 0</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,-153,228.5,-136</points>
<intersection>-153 3</intersection>
<intersection>-136 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>228,-136,228.5,-136</points>
<connection>
<GID>138</GID>
<name>OUT_1</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>228.5,-153,229.5,-153</points>
<connection>
<GID>137</GID>
<name>IN_1</name></connection>
<intersection>228.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-151,219,-134</points>
<connection>
<GID>140</GID>
<name>IN_3</name></connection>
<intersection>-147 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213.5,-147,219,-147</points>
<intersection>213.5 17</intersection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>217.5,-134,219,-134</points>
<connection>
<GID>141</GID>
<name>OUT_3</name></connection>
<intersection>219 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>213.5,-147,213.5,-146.5</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>-147 1</intersection></vsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217.5,-154,217.5,-137</points>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection>
<intersection>-154 5</intersection>
<intersection>-146.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>215.5,-146.5,217.5,-146.5</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>217.5,-154,219,-154</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-152,218.5,-135</points>
<intersection>-152 1</intersection>
<intersection>-135 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218.5,-152,219,-152</points>
<connection>
<GID>140</GID>
<name>IN_2</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>217.5,-135,218.5,-135</points>
<connection>
<GID>141</GID>
<name>OUT_2</name></connection>
<intersection>218.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-153,218,-136</points>
<intersection>-153 3</intersection>
<intersection>-136 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>217.5,-136,218,-136</points>
<connection>
<GID>141</GID>
<name>OUT_1</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>218,-153,219,-153</points>
<connection>
<GID>140</GID>
<name>IN_1</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209,-140,209,-130.5</points>
<intersection>-140 4</intersection>
<intersection>-130.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>209,-130.5,213.5,-130.5</points>
<intersection>209 0</intersection>
<intersection>213.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>209,-140,225,-140</points>
<connection>
<GID>141</GID>
<name>clock</name></connection>
<intersection>209 0</intersection>
<intersection>225 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>225,-140.5,225,-140</points>
<connection>
<GID>139</GID>
<name>OUT</name></connection>
<connection>
<GID>138</GID>
<name>clear</name></connection>
<intersection>-140 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>213.5,-131,213.5,-130.5</points>
<connection>
<GID>141</GID>
<name>count_enable</name></connection>
<intersection>-130.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-151,208.5,-134</points>
<connection>
<GID>143</GID>
<name>IN_3</name></connection>
<intersection>-147 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-147,208.5,-147</points>
<intersection>203 17</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207,-134,208.5,-134</points>
<connection>
<GID>144</GID>
<name>OUT_3</name></connection>
<intersection>208.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>203,-147,203,-146.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>-147 1</intersection></vsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-154,207,-137</points>
<connection>
<GID>144</GID>
<name>OUT_0</name></connection>
<intersection>-154 5</intersection>
<intersection>-146.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>205,-146.5,207,-146.5</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>207,-154,208.5,-154</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-152,208,-135</points>
<intersection>-152 1</intersection>
<intersection>-135 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208,-152,208.5,-152</points>
<connection>
<GID>143</GID>
<name>IN_2</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207,-135,208,-135</points>
<connection>
<GID>144</GID>
<name>OUT_2</name></connection>
<intersection>208 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,-153,207.5,-136</points>
<intersection>-153 3</intersection>
<intersection>-136 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>207,-136,207.5,-136</points>
<connection>
<GID>144</GID>
<name>OUT_1</name></connection>
<intersection>207.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>207.5,-153,208.5,-153</points>
<connection>
<GID>143</GID>
<name>IN_1</name></connection>
<intersection>207.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-140.5,198.5,-130.5</points>
<intersection>-140.5 4</intersection>
<intersection>-130.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198.5,-130.5,203,-130.5</points>
<intersection>198.5 0</intersection>
<intersection>203 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>198.5,-140.5,214.5,-140.5</points>
<intersection>198.5 0</intersection>
<intersection>202 15</intersection>
<intersection>214.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>214.5,-140.5,214.5,-140</points>
<connection>
<GID>142</GID>
<name>OUT</name></connection>
<connection>
<GID>141</GID>
<name>clear</name></connection>
<intersection>-140.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>203,-131,203,-130.5</points>
<connection>
<GID>144</GID>
<name>count_enable</name></connection>
<intersection>-130.5 3</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>202,-140.5,202,-140</points>
<connection>
<GID>144</GID>
<name>clock</name></connection>
<intersection>-140.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>256.5,-140.5,256.5,-140</points>
<connection>
<GID>130</GID>
<name>OUT</name></connection>
<connection>
<GID>129</GID>
<name>clear</name></connection>
<intersection>-140.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>240.5,-140.5,256.5,-140.5</points>
<intersection>240.5 4</intersection>
<intersection>244 8</intersection>
<intersection>256.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>240.5,-140.5,240.5,-130.5</points>
<intersection>-140.5 3</intersection>
<intersection>-130.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>240.5,-130.5,245,-130.5</points>
<intersection>240.5 4</intersection>
<intersection>245 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>245,-131,245,-130.5</points>
<connection>
<GID>132</GID>
<name>count_enable</name></connection>
<intersection>-130.5 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>244,-140.5,244,-140</points>
<connection>
<GID>132</GID>
<name>clock</name></connection>
<intersection>-140.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-140.5,246,-140</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<connection>
<GID>132</GID>
<name>clear</name></connection>
<intersection>-140.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230,-140.5,246,-140.5</points>
<intersection>230 4</intersection>
<intersection>233.5 20</intersection>
<intersection>246 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>230,-140.5,230,-131</points>
<intersection>-140.5 1</intersection>
<intersection>-131 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>230,-131,234.5,-131</points>
<connection>
<GID>135</GID>
<name>count_enable</name></connection>
<intersection>230 4</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>233.5,-140.5,233.5,-140</points>
<connection>
<GID>135</GID>
<name>clock</name></connection>
<intersection>-140.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303,-97,303,-80</points>
<connection>
<GID>146</GID>
<name>IN_3</name></connection>
<intersection>-93 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>297.5,-93,303,-93</points>
<intersection>297.5 17</intersection>
<intersection>303 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301.5,-80,303,-80</points>
<connection>
<GID>147</GID>
<name>OUT_3</name></connection>
<intersection>303 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>297.5,-93,297.5,-92.5</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-100,301.5,-83</points>
<connection>
<GID>147</GID>
<name>OUT_0</name></connection>
<intersection>-100 5</intersection>
<intersection>-92.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>299.5,-92.5,301.5,-92.5</points>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>301.5,-100,303,-100</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,-98,302.5,-81</points>
<intersection>-98 1</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302.5,-98,303,-98</points>
<connection>
<GID>146</GID>
<name>IN_2</name></connection>
<intersection>302.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301.5,-81,302.5,-81</points>
<connection>
<GID>147</GID>
<name>OUT_2</name></connection>
<intersection>302.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-99,302,-82</points>
<intersection>-99 3</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>301.5,-82,302,-82</points>
<connection>
<GID>147</GID>
<name>OUT_1</name></connection>
<intersection>302 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>302,-99,303,-99</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>302 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298.5,-86.5,298.5,-86</points>
<connection>
<GID>148</GID>
<name>OUT</name></connection>
<connection>
<GID>147</GID>
<name>clear</name></connection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282.5,-86.5,298.5,-86.5</points>
<intersection>282.5 2</intersection>
<intersection>286 7</intersection>
<intersection>298.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>282.5,-86.5,282.5,-76.5</points>
<intersection>-86.5 1</intersection>
<intersection>-76.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>282.5,-76.5,287,-76.5</points>
<intersection>282.5 2</intersection>
<intersection>287 10</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>286,-86.5,286,-86</points>
<connection>
<GID>150</GID>
<name>clock</name></connection>
<intersection>-86.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>287,-77,287,-76.5</points>
<connection>
<GID>150</GID>
<name>count_enable</name></connection>
<intersection>-76.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,-97,292.5,-80</points>
<connection>
<GID>149</GID>
<name>IN_3</name></connection>
<intersection>-93 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287,-93,292.5,-93</points>
<intersection>287 17</intersection>
<intersection>292.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>291,-80,292.5,-80</points>
<connection>
<GID>150</GID>
<name>OUT_3</name></connection>
<intersection>292.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>287,-93,287,-92.5</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,-100,291,-83</points>
<connection>
<GID>150</GID>
<name>OUT_0</name></connection>
<intersection>-100 5</intersection>
<intersection>-92.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>289,-92.5,291,-92.5</points>
<connection>
<GID>151</GID>
<name>IN_1</name></connection>
<intersection>291 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>291,-100,292.5,-100</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>291 0</intersection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,-98,292,-81</points>
<intersection>-98 1</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>292,-98,292.5,-98</points>
<connection>
<GID>149</GID>
<name>IN_2</name></connection>
<intersection>292 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>291,-81,292,-81</points>
<connection>
<GID>150</GID>
<name>OUT_2</name></connection>
<intersection>292 0</intersection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,-99,291.5,-82</points>
<intersection>-99 3</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>291,-82,291.5,-82</points>
<connection>
<GID>150</GID>
<name>OUT_1</name></connection>
<intersection>291.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>291.5,-99,292.5,-99</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,-86.5,288,-86</points>
<connection>
<GID>151</GID>
<name>OUT</name></connection>
<connection>
<GID>150</GID>
<name>clear</name></connection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>272,-86.5,288,-86.5</points>
<intersection>272 2</intersection>
<intersection>275.5 12</intersection>
<intersection>288 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>272,-86.5,272,-77</points>
<intersection>-86.5 1</intersection>
<intersection>-77 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>272,-77,276.5,-77</points>
<connection>
<GID>153</GID>
<name>count_enable</name></connection>
<intersection>272 2</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>275.5,-86.5,275.5,-86</points>
<connection>
<GID>153</GID>
<name>clock</name></connection>
<intersection>-86.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-97,282,-80</points>
<connection>
<GID>152</GID>
<name>IN_3</name></connection>
<intersection>-93 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276.5,-93,282,-93</points>
<intersection>276.5 17</intersection>
<intersection>282 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280.5,-80,282,-80</points>
<connection>
<GID>153</GID>
<name>OUT_3</name></connection>
<intersection>282 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>276.5,-93,276.5,-92.5</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280.5,-100,280.5,-83</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>-100 5</intersection>
<intersection>-92.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>278.5,-92.5,280.5,-92.5</points>
<connection>
<GID>154</GID>
<name>IN_1</name></connection>
<intersection>280.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>280.5,-100,282,-100</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>280.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-98,281.5,-81</points>
<intersection>-98 1</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281.5,-98,282,-98</points>
<connection>
<GID>152</GID>
<name>IN_2</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280.5,-81,281.5,-81</points>
<connection>
<GID>153</GID>
<name>OUT_2</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,-99,281,-82</points>
<intersection>-99 3</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>280.5,-82,281,-82</points>
<connection>
<GID>153</GID>
<name>OUT_1</name></connection>
<intersection>281 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>281,-99,282,-99</points>
<connection>
<GID>152</GID>
<name>IN_1</name></connection>
<intersection>281 0</intersection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,-97,271.5,-80</points>
<connection>
<GID>155</GID>
<name>IN_3</name></connection>
<intersection>-93 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266,-93,271.5,-93</points>
<intersection>266 17</intersection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>270,-80,271.5,-80</points>
<connection>
<GID>186</GID>
<name>OUT_3</name></connection>
<intersection>271.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>266,-93,266,-92.5</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,-100,270,-83</points>
<connection>
<GID>186</GID>
<name>OUT_0</name></connection>
<intersection>-100 5</intersection>
<intersection>-92.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>268,-92.5,270,-92.5</points>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<intersection>270 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>270,-100,271.5,-100</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>270 0</intersection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-98,271,-81</points>
<intersection>-98 1</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>271,-98,271.5,-98</points>
<connection>
<GID>155</GID>
<name>IN_2</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>270,-81,271,-81</points>
<connection>
<GID>186</GID>
<name>OUT_2</name></connection>
<intersection>271 0</intersection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-99,270.5,-82</points>
<intersection>-99 3</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>270,-82,270.5,-82</points>
<connection>
<GID>186</GID>
<name>OUT_1</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>270.5,-99,271.5,-99</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,-86.5,261.5,-76.5</points>
<intersection>-86.5 4</intersection>
<intersection>-76.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>261.5,-76.5,266,-76.5</points>
<intersection>261.5 0</intersection>
<intersection>266 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>261.5,-86.5,277.5,-86.5</points>
<intersection>261.5 0</intersection>
<intersection>265 7</intersection>
<intersection>277.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>277.5,-86.5,277.5,-86</points>
<connection>
<GID>154</GID>
<name>OUT</name></connection>
<connection>
<GID>153</GID>
<name>clear</name></connection>
<intersection>-86.5 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>265,-86.5,265,-86</points>
<connection>
<GID>186</GID>
<name>clock</name></connection>
<intersection>-86.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>266,-77,266,-76.5</points>
<connection>
<GID>186</GID>
<name>count_enable</name></connection>
<intersection>-76.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,-97,261,-80</points>
<connection>
<GID>188</GID>
<name>IN_3</name></connection>
<intersection>-93 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255.5,-93,261,-93</points>
<intersection>255.5 17</intersection>
<intersection>261 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259.5,-80,261,-80</points>
<connection>
<GID>189</GID>
<name>OUT_3</name></connection>
<intersection>261 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>255.5,-93,255.5,-92.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,-100,259.5,-83</points>
<connection>
<GID>189</GID>
<name>OUT_0</name></connection>
<intersection>-100 5</intersection>
<intersection>-92.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>257.5,-92.5,259.5,-92.5</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>259.5,-100,261,-100</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>259.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,-98,260.5,-81</points>
<intersection>-98 1</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,-98,261,-98</points>
<connection>
<GID>188</GID>
<name>IN_2</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259.5,-81,260.5,-81</points>
<connection>
<GID>189</GID>
<name>OUT_2</name></connection>
<intersection>260.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-99,260,-82</points>
<intersection>-99 3</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>259.5,-82,260,-82</points>
<connection>
<GID>189</GID>
<name>OUT_1</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>260,-99,261,-99</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,-86,251,-76.5</points>
<intersection>-86 4</intersection>
<intersection>-76.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>251,-76.5,255.5,-76.5</points>
<intersection>251 0</intersection>
<intersection>255.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>251,-86,267,-86</points>
<connection>
<GID>189</GID>
<name>clock</name></connection>
<intersection>251 0</intersection>
<intersection>267 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>267,-86.5,267,-86</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<connection>
<GID>186</GID>
<name>clear</name></connection>
<intersection>-86 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>255.5,-77,255.5,-76.5</points>
<connection>
<GID>189</GID>
<name>count_enable</name></connection>
<intersection>-76.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-86,293,-76.5</points>
<intersection>-86 4</intersection>
<intersection>-76.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>293,-76.5,297.5,-76.5</points>
<intersection>293 0</intersection>
<intersection>297.5 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293,-86,296.5,-86</points>
<connection>
<GID>147</GID>
<name>clock</name></connection>
<intersection>293 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>297.5,-77,297.5,-76</points>
<connection>
<GID>147</GID>
<name>count_enable</name></connection>
<intersection>-76.5 3</intersection>
<intersection>-76 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>197.5,-76,297.5,-76</points>
<intersection>197.5 7</intersection>
<intersection>297.5 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>197.5,-113.5,197.5,-76</points>
<intersection>-113.5 8</intersection>
<intersection>-76 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>197.5,-113.5,204,-113.5</points>
<connection>
<GID>124</GID>
<name>clear</name></connection>
<intersection>197.5 7</intersection>
<intersection>204 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>204,-114,204,-113.5</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>-113.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,-97,250.5,-80</points>
<connection>
<GID>191</GID>
<name>IN_3</name></connection>
<intersection>-93 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245,-93,250.5,-93</points>
<intersection>245 17</intersection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>249,-80,250.5,-80</points>
<connection>
<GID>192</GID>
<name>OUT_3</name></connection>
<intersection>250.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>245,-93,245,-92.5</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303,-70.5,303,-53.5</points>
<connection>
<GID>156</GID>
<name>IN_3</name></connection>
<intersection>-66.5 1</intersection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>297.5,-66.5,303,-66.5</points>
<intersection>297.5 17</intersection>
<intersection>303 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301.5,-53.5,303,-53.5</points>
<connection>
<GID>157</GID>
<name>OUT_3</name></connection>
<intersection>303 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>297.5,-66.5,297.5,-66</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>-66.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-73.5,301.5,-56.5</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>-73.5 5</intersection>
<intersection>-66 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>299.5,-66,301.5,-66</points>
<connection>
<GID>158</GID>
<name>IN_1</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>301.5,-73.5,303,-73.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,-71.5,302.5,-54.5</points>
<intersection>-71.5 1</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302.5,-71.5,303,-71.5</points>
<connection>
<GID>156</GID>
<name>IN_2</name></connection>
<intersection>302.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301.5,-54.5,302.5,-54.5</points>
<connection>
<GID>157</GID>
<name>OUT_2</name></connection>
<intersection>302.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-72.5,302,-55.5</points>
<intersection>-72.5 3</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>301.5,-55.5,302,-55.5</points>
<connection>
<GID>157</GID>
<name>OUT_1</name></connection>
<intersection>302 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>302,-72.5,303,-72.5</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<intersection>302 0</intersection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298.5,-60,298.5,-59.5</points>
<connection>
<GID>158</GID>
<name>OUT</name></connection>
<connection>
<GID>157</GID>
<name>clear</name></connection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282.5,-60,298.5,-60</points>
<intersection>282.5 2</intersection>
<intersection>286 7</intersection>
<intersection>298.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>282.5,-60,282.5,-50</points>
<intersection>-60 1</intersection>
<intersection>-50 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>282.5,-50,287,-50</points>
<intersection>282.5 2</intersection>
<intersection>287 10</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>286,-60,286,-59.5</points>
<connection>
<GID>160</GID>
<name>clock</name></connection>
<intersection>-60 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>287,-50.5,287,-50</points>
<connection>
<GID>160</GID>
<name>count_enable</name></connection>
<intersection>-50 5</intersection></vsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249,-100,249,-83</points>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection>
<intersection>-100 5</intersection>
<intersection>-92.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>247,-92.5,249,-92.5</points>
<connection>
<GID>193</GID>
<name>IN_1</name></connection>
<intersection>249 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>249,-100,250.5,-100</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>249 0</intersection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,-70.5,292.5,-53.5</points>
<connection>
<GID>159</GID>
<name>IN_3</name></connection>
<intersection>-66.5 1</intersection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287,-66.5,292.5,-66.5</points>
<intersection>287 17</intersection>
<intersection>292.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>291,-53.5,292.5,-53.5</points>
<connection>
<GID>160</GID>
<name>OUT_3</name></connection>
<intersection>292.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>287,-66.5,287,-66</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>-66.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,-73.5,291,-56.5</points>
<connection>
<GID>160</GID>
<name>OUT_0</name></connection>
<intersection>-73.5 5</intersection>
<intersection>-66 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>289,-66,291,-66</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<intersection>291 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>291,-73.5,292.5,-73.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>291 0</intersection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,-71.5,292,-54.5</points>
<intersection>-71.5 1</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>292,-71.5,292.5,-71.5</points>
<connection>
<GID>159</GID>
<name>IN_2</name></connection>
<intersection>292 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>291,-54.5,292,-54.5</points>
<connection>
<GID>160</GID>
<name>OUT_2</name></connection>
<intersection>292 0</intersection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,-72.5,291.5,-55.5</points>
<intersection>-72.5 3</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>291,-55.5,291.5,-55.5</points>
<connection>
<GID>160</GID>
<name>OUT_1</name></connection>
<intersection>291.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>291.5,-72.5,292.5,-72.5</points>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,-60,288,-59.5</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<connection>
<GID>160</GID>
<name>clear</name></connection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>272,-59.5,288,-59.5</points>
<connection>
<GID>163</GID>
<name>clock</name></connection>
<intersection>272 2</intersection>
<intersection>288 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>272,-59.5,272,-50</points>
<intersection>-59.5 1</intersection>
<intersection>-50 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>272,-50,276.5,-50</points>
<intersection>272 2</intersection>
<intersection>276.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>276.5,-50.5,276.5,-50</points>
<connection>
<GID>163</GID>
<name>count_enable</name></connection>
<intersection>-50 5</intersection></vsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-70.5,282,-53.5</points>
<connection>
<GID>162</GID>
<name>IN_3</name></connection>
<intersection>-66.5 1</intersection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276.5,-66.5,282,-66.5</points>
<intersection>276.5 17</intersection>
<intersection>282 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280.5,-53.5,282,-53.5</points>
<connection>
<GID>163</GID>
<name>OUT_3</name></connection>
<intersection>282 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>276.5,-66.5,276.5,-66</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>-66.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280.5,-73.5,280.5,-56.5</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>-73.5 5</intersection>
<intersection>-66 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>278.5,-66,280.5,-66</points>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<intersection>280.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>280.5,-73.5,282,-73.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>280.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-71.5,281.5,-54.5</points>
<intersection>-71.5 1</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281.5,-71.5,282,-71.5</points>
<connection>
<GID>162</GID>
<name>IN_2</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280.5,-54.5,281.5,-54.5</points>
<connection>
<GID>163</GID>
<name>OUT_2</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,-72.5,281,-55.5</points>
<intersection>-72.5 3</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>280.5,-55.5,281,-55.5</points>
<connection>
<GID>163</GID>
<name>OUT_1</name></connection>
<intersection>281 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>281,-72.5,282,-72.5</points>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<intersection>281 0</intersection></hsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,-70.5,271.5,-53.5</points>
<connection>
<GID>165</GID>
<name>IN_3</name></connection>
<intersection>-66.5 1</intersection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266,-66.5,271.5,-66.5</points>
<intersection>266 17</intersection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>270,-53.5,271.5,-53.5</points>
<connection>
<GID>166</GID>
<name>OUT_3</name></connection>
<intersection>271.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>266,-66.5,266,-66</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>-66.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,-73.5,270,-56.5</points>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection>
<intersection>-73.5 5</intersection>
<intersection>-66 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>268,-66,270,-66</points>
<connection>
<GID>167</GID>
<name>IN_1</name></connection>
<intersection>270 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>270,-73.5,271.5,-73.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>270 0</intersection></hsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-71.5,271,-54.5</points>
<intersection>-71.5 1</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>271,-71.5,271.5,-71.5</points>
<connection>
<GID>165</GID>
<name>IN_2</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>270,-54.5,271,-54.5</points>
<connection>
<GID>166</GID>
<name>OUT_2</name></connection>
<intersection>271 0</intersection></hsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-72.5,270.5,-55.5</points>
<intersection>-72.5 3</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>270,-55.5,270.5,-55.5</points>
<connection>
<GID>166</GID>
<name>OUT_1</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>270.5,-72.5,271.5,-72.5</points>
<connection>
<GID>165</GID>
<name>IN_1</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,-60,261.5,-50</points>
<intersection>-60 4</intersection>
<intersection>-50 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>261.5,-50,266,-50</points>
<intersection>261.5 0</intersection>
<intersection>266 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>261.5,-60,277.5,-60</points>
<intersection>261.5 0</intersection>
<intersection>265 7</intersection>
<intersection>277.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>277.5,-60,277.5,-59.5</points>
<connection>
<GID>164</GID>
<name>OUT</name></connection>
<connection>
<GID>163</GID>
<name>clear</name></connection>
<intersection>-60 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>265,-60,265,-59.5</points>
<connection>
<GID>166</GID>
<name>clock</name></connection>
<intersection>-60 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>266,-50.5,266,-50</points>
<connection>
<GID>166</GID>
<name>count_enable</name></connection>
<intersection>-50 3</intersection></vsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,-70.5,261,-53.5</points>
<connection>
<GID>168</GID>
<name>IN_3</name></connection>
<intersection>-66.5 1</intersection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255.5,-66.5,261,-66.5</points>
<intersection>255.5 17</intersection>
<intersection>261 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259.5,-53.5,261,-53.5</points>
<connection>
<GID>169</GID>
<name>OUT_3</name></connection>
<intersection>261 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>255.5,-66.5,255.5,-66</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>-66.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,-73.5,259.5,-56.5</points>
<connection>
<GID>169</GID>
<name>OUT_0</name></connection>
<intersection>-73.5 5</intersection>
<intersection>-66 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>257.5,-66,259.5,-66</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>259.5,-73.5,261,-73.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>259.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,-71.5,260.5,-54.5</points>
<intersection>-71.5 1</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,-71.5,261,-71.5</points>
<connection>
<GID>168</GID>
<name>IN_2</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259.5,-54.5,260.5,-54.5</points>
<connection>
<GID>169</GID>
<name>OUT_2</name></connection>
<intersection>260.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-72.5,260,-55.5</points>
<intersection>-72.5 3</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>259.5,-55.5,260,-55.5</points>
<connection>
<GID>169</GID>
<name>OUT_1</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>260,-72.5,261,-72.5</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,-98,250,-81</points>
<intersection>-98 1</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250,-98,250.5,-98</points>
<connection>
<GID>191</GID>
<name>IN_2</name></connection>
<intersection>250 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>249,-81,250,-81</points>
<connection>
<GID>192</GID>
<name>OUT_2</name></connection>
<intersection>250 0</intersection></hsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,-59.5,251,-50</points>
<intersection>-59.5 4</intersection>
<intersection>-50 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>251,-50,255.5,-50</points>
<intersection>251 0</intersection>
<intersection>255.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>251,-59.5,267,-59.5</points>
<connection>
<GID>169</GID>
<name>clock</name></connection>
<intersection>251 0</intersection>
<intersection>267 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>267,-60,267,-59.5</points>
<connection>
<GID>167</GID>
<name>OUT</name></connection>
<connection>
<GID>166</GID>
<name>clear</name></connection>
<intersection>-59.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>255.5,-50.5,255.5,-50</points>
<connection>
<GID>169</GID>
<name>count_enable</name></connection>
<intersection>-50 3</intersection></vsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-59.5,293,-50</points>
<intersection>-59.5 4</intersection>
<intersection>-50 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>293,-50,297.5,-50</points>
<intersection>293 0</intersection>
<intersection>297.5 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293,-59.5,296.5,-59.5</points>
<connection>
<GID>157</GID>
<name>clock</name></connection>
<intersection>293 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>297.5,-50.5,297.5,-49</points>
<connection>
<GID>157</GID>
<name>count_enable</name></connection>
<intersection>-50 3</intersection>
<intersection>-49 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>196.5,-49,297.5,-49</points>
<intersection>196.5 7</intersection>
<intersection>297.5 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>196.5,-86.5,196.5,-49</points>
<intersection>-86.5 8</intersection>
<intersection>-49 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>196.5,-86.5,204,-86.5</points>
<connection>
<GID>205</GID>
<name>OUT</name></connection>
<intersection>196.5 7</intersection>
<intersection>204 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>204,-86.5,204,-86</points>
<connection>
<GID>204</GID>
<name>clear</name></connection>
<intersection>-86.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,-70.5,250.5,-53.5</points>
<connection>
<GID>171</GID>
<name>IN_3</name></connection>
<intersection>-66.5 1</intersection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245,-66.5,250.5,-66.5</points>
<intersection>245 17</intersection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>249,-53.5,250.5,-53.5</points>
<connection>
<GID>172</GID>
<name>OUT_3</name></connection>
<intersection>250.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>245,-66.5,245,-66</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>-66.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249,-73.5,249,-56.5</points>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection>
<intersection>-73.5 5</intersection>
<intersection>-66 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>247,-66,249,-66</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<intersection>249 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>249,-73.5,250.5,-73.5</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>249 0</intersection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,-71.5,250,-54.5</points>
<intersection>-71.5 1</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250,-71.5,250.5,-71.5</points>
<connection>
<GID>171</GID>
<name>IN_2</name></connection>
<intersection>250 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>249,-54.5,250,-54.5</points>
<connection>
<GID>172</GID>
<name>OUT_2</name></connection>
<intersection>250 0</intersection></hsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,-72.5,249.5,-55.5</points>
<intersection>-72.5 3</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>249,-55.5,249.5,-55.5</points>
<connection>
<GID>172</GID>
<name>OUT_1</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>249.5,-72.5,250.5,-72.5</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<intersection>249.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,-99,249.5,-82</points>
<intersection>-99 3</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>249,-82,249.5,-82</points>
<connection>
<GID>192</GID>
<name>OUT_1</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>249.5,-99,250.5,-99</points>
<connection>
<GID>191</GID>
<name>IN_1</name></connection>
<intersection>249.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-70.5,240,-53.5</points>
<connection>
<GID>174</GID>
<name>IN_3</name></connection>
<intersection>-66.5 1</intersection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234.5,-66.5,240,-66.5</points>
<intersection>234.5 17</intersection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-53.5,240,-53.5</points>
<connection>
<GID>175</GID>
<name>OUT_3</name></connection>
<intersection>240 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>234.5,-66.5,234.5,-66</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>-66.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,-73.5,238.5,-56.5</points>
<connection>
<GID>175</GID>
<name>OUT_0</name></connection>
<intersection>-73.5 5</intersection>
<intersection>-66 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>236.5,-66,238.5,-66</points>
<connection>
<GID>176</GID>
<name>IN_1</name></connection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>238.5,-73.5,240,-73.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>238.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239.5,-71.5,239.5,-54.5</points>
<intersection>-71.5 1</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239.5,-71.5,240,-71.5</points>
<connection>
<GID>174</GID>
<name>IN_2</name></connection>
<intersection>239.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-54.5,239.5,-54.5</points>
<connection>
<GID>175</GID>
<name>OUT_2</name></connection>
<intersection>239.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,-72.5,239,-55.5</points>
<intersection>-72.5 3</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-55.5,239,-55.5</points>
<connection>
<GID>175</GID>
<name>OUT_1</name></connection>
<intersection>239 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>239,-72.5,240,-72.5</points>
<connection>
<GID>174</GID>
<name>IN_1</name></connection>
<intersection>239 0</intersection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235.5,-60,235.5,-59.5</points>
<connection>
<GID>176</GID>
<name>OUT</name></connection>
<connection>
<GID>175</GID>
<name>clear</name></connection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219.5,-60,235.5,-60</points>
<intersection>219.5 2</intersection>
<intersection>223 10</intersection>
<intersection>235.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>219.5,-60,219.5,-50</points>
<intersection>-60 1</intersection>
<intersection>-50 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>219.5,-50,224,-50</points>
<intersection>219.5 2</intersection>
<intersection>224 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>224,-50.5,224,-50</points>
<connection>
<GID>178</GID>
<name>count_enable</name></connection>
<intersection>-50 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>223,-60,223,-59.5</points>
<connection>
<GID>178</GID>
<name>clock</name></connection>
<intersection>-60 1</intersection></vsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,-70.5,229.5,-53.5</points>
<connection>
<GID>177</GID>
<name>IN_3</name></connection>
<intersection>-66.5 1</intersection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>224,-66.5,229.5,-66.5</points>
<intersection>224 17</intersection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228,-53.5,229.5,-53.5</points>
<connection>
<GID>178</GID>
<name>OUT_3</name></connection>
<intersection>229.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>224,-66.5,224,-66</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>-66.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,-73.5,228,-56.5</points>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<intersection>-73.5 5</intersection>
<intersection>-66 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-66,228,-66</points>
<connection>
<GID>179</GID>
<name>IN_1</name></connection>
<intersection>228 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>228,-73.5,229.5,-73.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>228 0</intersection></hsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-71.5,229,-54.5</points>
<intersection>-71.5 1</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229,-71.5,229.5,-71.5</points>
<connection>
<GID>177</GID>
<name>IN_2</name></connection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228,-54.5,229,-54.5</points>
<connection>
<GID>178</GID>
<name>OUT_2</name></connection>
<intersection>229 0</intersection></hsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,-72.5,228.5,-55.5</points>
<intersection>-72.5 3</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>228,-55.5,228.5,-55.5</points>
<connection>
<GID>178</GID>
<name>OUT_1</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>228.5,-72.5,229.5,-72.5</points>
<connection>
<GID>177</GID>
<name>IN_1</name></connection>
<intersection>228.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-70.5,219,-53.5</points>
<connection>
<GID>180</GID>
<name>IN_3</name></connection>
<intersection>-66.5 1</intersection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213.5,-66.5,219,-66.5</points>
<intersection>213.5 17</intersection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>217.5,-53.5,219,-53.5</points>
<connection>
<GID>181</GID>
<name>OUT_3</name></connection>
<intersection>219 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>213.5,-66.5,213.5,-66</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>-66.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217.5,-73.5,217.5,-56.5</points>
<connection>
<GID>181</GID>
<name>OUT_0</name></connection>
<intersection>-73.5 5</intersection>
<intersection>-66 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>215.5,-66,217.5,-66</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>217.5,-73.5,219,-73.5</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-71.5,218.5,-54.5</points>
<intersection>-71.5 1</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218.5,-71.5,219,-71.5</points>
<connection>
<GID>180</GID>
<name>IN_2</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>217.5,-54.5,218.5,-54.5</points>
<connection>
<GID>181</GID>
<name>OUT_2</name></connection>
<intersection>218.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-72.5,218,-55.5</points>
<intersection>-72.5 3</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>217.5,-55.5,218,-55.5</points>
<connection>
<GID>181</GID>
<name>OUT_1</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>218,-72.5,219,-72.5</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209,-59.5,209,-50</points>
<intersection>-59.5 4</intersection>
<intersection>-50 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>209,-50,213.5,-50</points>
<intersection>209 0</intersection>
<intersection>213.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>209,-59.5,225,-59.5</points>
<connection>
<GID>181</GID>
<name>clock</name></connection>
<intersection>209 0</intersection>
<intersection>225 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>225,-60,225,-59.5</points>
<connection>
<GID>179</GID>
<name>OUT</name></connection>
<connection>
<GID>178</GID>
<name>clear</name></connection>
<intersection>-59.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>213.5,-50.5,213.5,-50</points>
<connection>
<GID>181</GID>
<name>count_enable</name></connection>
<intersection>-50 3</intersection></vsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-70.5,208.5,-53.5</points>
<connection>
<GID>183</GID>
<name>IN_3</name></connection>
<intersection>-66.5 1</intersection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-66.5,208.5,-66.5</points>
<intersection>203 17</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207,-53.5,208.5,-53.5</points>
<connection>
<GID>184</GID>
<name>OUT_3</name></connection>
<intersection>208.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>203,-66.5,203,-66</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>-66.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-73.5,207,-56.5</points>
<connection>
<GID>184</GID>
<name>OUT_0</name></connection>
<intersection>-73.5 5</intersection>
<intersection>-66 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>205,-66,207,-66</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>207,-73.5,208.5,-73.5</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-71.5,208,-54.5</points>
<intersection>-71.5 1</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208,-71.5,208.5,-71.5</points>
<connection>
<GID>183</GID>
<name>IN_2</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207,-54.5,208,-54.5</points>
<connection>
<GID>184</GID>
<name>OUT_2</name></connection>
<intersection>208 0</intersection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,-72.5,207.5,-55.5</points>
<intersection>-72.5 3</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>207,-55.5,207.5,-55.5</points>
<connection>
<GID>184</GID>
<name>OUT_1</name></connection>
<intersection>207.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>207.5,-72.5,208.5,-72.5</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>207.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-60,198.5,-50</points>
<intersection>-60 4</intersection>
<intersection>-50 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198.5,-50,203,-50</points>
<intersection>198.5 0</intersection>
<intersection>203 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>198.5,-60,214.5,-60</points>
<intersection>198.5 0</intersection>
<intersection>202 15</intersection>
<intersection>214.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>214.5,-60,214.5,-59.5</points>
<connection>
<GID>182</GID>
<name>OUT</name></connection>
<connection>
<GID>181</GID>
<name>clear</name></connection>
<intersection>-60 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>203,-50.5,203,-50</points>
<connection>
<GID>184</GID>
<name>count_enable</name></connection>
<intersection>-50 3</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>202,-60,202,-59.5</points>
<connection>
<GID>184</GID>
<name>clock</name></connection>
<intersection>-60 4</intersection></vsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-97,240,-80</points>
<connection>
<GID>194</GID>
<name>IN_3</name></connection>
<intersection>-93 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234.5,-93,240,-93</points>
<intersection>234.5 17</intersection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-80,240,-80</points>
<connection>
<GID>195</GID>
<name>OUT_3</name></connection>
<intersection>240 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>234.5,-93,234.5,-92.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>256.5,-60,256.5,-59.5</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<connection>
<GID>169</GID>
<name>clear</name></connection>
<intersection>-60 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>240.5,-60,256.5,-60</points>
<intersection>240.5 4</intersection>
<intersection>244 8</intersection>
<intersection>256.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>240.5,-60,240.5,-50</points>
<intersection>-60 3</intersection>
<intersection>-50 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>240.5,-50,245,-50</points>
<intersection>240.5 4</intersection>
<intersection>245 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>245,-50.5,245,-50</points>
<connection>
<GID>172</GID>
<name>count_enable</name></connection>
<intersection>-50 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>244,-60,244,-59.5</points>
<connection>
<GID>172</GID>
<name>clock</name></connection>
<intersection>-60 3</intersection></vsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-60,246,-59.5</points>
<connection>
<GID>173</GID>
<name>OUT</name></connection>
<connection>
<GID>172</GID>
<name>clear</name></connection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230,-59.5,246,-59.5</points>
<connection>
<GID>175</GID>
<name>clock</name></connection>
<intersection>230 4</intersection>
<intersection>246 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>230,-59.5,230,-50</points>
<intersection>-59.5 1</intersection>
<intersection>-50 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>230,-50,234.5,-50</points>
<intersection>230 4</intersection>
<intersection>234.5 17</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>234.5,-50.5,234.5,-50</points>
<connection>
<GID>175</GID>
<name>count_enable</name></connection>
<intersection>-50 15</intersection></vsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,-100,238.5,-83</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<intersection>-100 5</intersection>
<intersection>-92.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>236.5,-92.5,238.5,-92.5</points>
<connection>
<GID>196</GID>
<name>IN_1</name></connection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>238.5,-100,240,-100</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>238.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239.5,-98,239.5,-81</points>
<intersection>-98 1</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239.5,-98,240,-98</points>
<connection>
<GID>194</GID>
<name>IN_2</name></connection>
<intersection>239.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-81,239.5,-81</points>
<connection>
<GID>195</GID>
<name>OUT_2</name></connection>
<intersection>239.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,-99,239,-82</points>
<intersection>-99 3</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-82,239,-82</points>
<connection>
<GID>195</GID>
<name>OUT_1</name></connection>
<intersection>239 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>239,-99,240,-99</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<intersection>239 0</intersection></hsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235.5,-86.5,235.5,-86</points>
<connection>
<GID>196</GID>
<name>OUT</name></connection>
<connection>
<GID>195</GID>
<name>clear</name></connection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219.5,-86.5,235.5,-86.5</points>
<intersection>219.5 2</intersection>
<intersection>223 10</intersection>
<intersection>235.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>219.5,-86.5,219.5,-76.5</points>
<intersection>-86.5 1</intersection>
<intersection>-76.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>219.5,-76.5,224,-76.5</points>
<intersection>219.5 2</intersection>
<intersection>224 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>224,-77,224,-76.5</points>
<connection>
<GID>198</GID>
<name>count_enable</name></connection>
<intersection>-76.5 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>223,-86.5,223,-86</points>
<connection>
<GID>198</GID>
<name>clock</name></connection>
<intersection>-86.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,-97,229.5,-80</points>
<connection>
<GID>197</GID>
<name>IN_3</name></connection>
<intersection>-93 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>224,-93,229.5,-93</points>
<intersection>224 17</intersection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228,-80,229.5,-80</points>
<connection>
<GID>198</GID>
<name>OUT_3</name></connection>
<intersection>229.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>224,-93,224,-92.5</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,-100,228,-83</points>
<connection>
<GID>198</GID>
<name>OUT_0</name></connection>
<intersection>-100 5</intersection>
<intersection>-92.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-92.5,228,-92.5</points>
<connection>
<GID>199</GID>
<name>IN_1</name></connection>
<intersection>228 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>228,-100,229.5,-100</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>228 0</intersection></hsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-98,229,-81</points>
<intersection>-98 1</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229,-98,229.5,-98</points>
<connection>
<GID>197</GID>
<name>IN_2</name></connection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228,-81,229,-81</points>
<connection>
<GID>198</GID>
<name>OUT_2</name></connection>
<intersection>229 0</intersection></hsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,-99,228.5,-82</points>
<intersection>-99 3</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>228,-82,228.5,-82</points>
<connection>
<GID>198</GID>
<name>OUT_1</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>228.5,-99,229.5,-99</points>
<connection>
<GID>197</GID>
<name>IN_1</name></connection>
<intersection>228.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-97,219,-80</points>
<connection>
<GID>200</GID>
<name>IN_3</name></connection>
<intersection>-93 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213.5,-93,219,-93</points>
<intersection>213.5 17</intersection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>217.5,-80,219,-80</points>
<connection>
<GID>201</GID>
<name>OUT_3</name></connection>
<intersection>219 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>213.5,-93,213.5,-92.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217.5,-100,217.5,-83</points>
<connection>
<GID>201</GID>
<name>OUT_0</name></connection>
<intersection>-100 5</intersection>
<intersection>-92.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>215.5,-92.5,217.5,-92.5</points>
<connection>
<GID>202</GID>
<name>IN_1</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>217.5,-100,219,-100</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-98,218.5,-81</points>
<intersection>-98 1</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218.5,-98,219,-98</points>
<connection>
<GID>200</GID>
<name>IN_2</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>217.5,-81,218.5,-81</points>
<connection>
<GID>201</GID>
<name>OUT_2</name></connection>
<intersection>218.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-99,218,-82</points>
<intersection>-99 3</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>217.5,-82,218,-82</points>
<connection>
<GID>201</GID>
<name>OUT_1</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>218,-99,219,-99</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209,-86,209,-76.5</points>
<intersection>-86 4</intersection>
<intersection>-76.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>209,-76.5,213.5,-76.5</points>
<intersection>209 0</intersection>
<intersection>213.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>209,-86,225,-86</points>
<connection>
<GID>201</GID>
<name>clock</name></connection>
<intersection>209 0</intersection>
<intersection>225 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>225,-86.5,225,-86</points>
<connection>
<GID>199</GID>
<name>OUT</name></connection>
<connection>
<GID>198</GID>
<name>clear</name></connection>
<intersection>-86 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>213.5,-77,213.5,-76.5</points>
<connection>
<GID>201</GID>
<name>count_enable</name></connection>
<intersection>-76.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-97,208.5,-80</points>
<connection>
<GID>203</GID>
<name>IN_3</name></connection>
<intersection>-93 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-93,208.5,-93</points>
<intersection>203 17</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207,-80,208.5,-80</points>
<connection>
<GID>204</GID>
<name>OUT_3</name></connection>
<intersection>208.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>203,-93,203,-92.5</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-100,207,-83</points>
<connection>
<GID>204</GID>
<name>OUT_0</name></connection>
<intersection>-100 5</intersection>
<intersection>-92.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>205,-92.5,207,-92.5</points>
<connection>
<GID>205</GID>
<name>IN_1</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>207,-100,208.5,-100</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-98,208,-81</points>
<intersection>-98 1</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208,-98,208.5,-98</points>
<connection>
<GID>203</GID>
<name>IN_2</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207,-81,208,-81</points>
<connection>
<GID>204</GID>
<name>OUT_2</name></connection>
<intersection>208 0</intersection></hsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,-99,207.5,-82</points>
<intersection>-99 3</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>207,-82,207.5,-82</points>
<connection>
<GID>204</GID>
<name>OUT_1</name></connection>
<intersection>207.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>207.5,-99,208.5,-99</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<intersection>207.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-86.5,198.5,-76.5</points>
<intersection>-86.5 4</intersection>
<intersection>-76.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198.5,-76.5,203,-76.5</points>
<intersection>198.5 0</intersection>
<intersection>203 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>198.5,-86.5,214.5,-86.5</points>
<intersection>198.5 0</intersection>
<intersection>202 15</intersection>
<intersection>214.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>214.5,-86.5,214.5,-86</points>
<connection>
<GID>202</GID>
<name>OUT</name></connection>
<connection>
<GID>201</GID>
<name>clear</name></connection>
<intersection>-86.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>203,-77,203,-76.5</points>
<connection>
<GID>204</GID>
<name>count_enable</name></connection>
<intersection>-76.5 3</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>202,-86.5,202,-86</points>
<connection>
<GID>204</GID>
<name>clock</name></connection>
<intersection>-86.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>256.5,-86.5,256.5,-86</points>
<connection>
<GID>190</GID>
<name>OUT</name></connection>
<connection>
<GID>189</GID>
<name>clear</name></connection>
<intersection>-86.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>240.5,-86.5,256.5,-86.5</points>
<intersection>240.5 4</intersection>
<intersection>244 8</intersection>
<intersection>256.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>240.5,-86.5,240.5,-76.5</points>
<intersection>-86.5 3</intersection>
<intersection>-76.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>240.5,-76.5,245,-76.5</points>
<intersection>240.5 4</intersection>
<intersection>245 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>245,-77,245,-76.5</points>
<connection>
<GID>192</GID>
<name>count_enable</name></connection>
<intersection>-76.5 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>244,-86.5,244,-86</points>
<connection>
<GID>192</GID>
<name>clock</name></connection>
<intersection>-86.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-86.5,246,-86</points>
<connection>
<GID>193</GID>
<name>OUT</name></connection>
<connection>
<GID>192</GID>
<name>clear</name></connection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230,-86.5,246,-86.5</points>
<intersection>230 4</intersection>
<intersection>233.5 20</intersection>
<intersection>246 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>230,-86.5,230,-77</points>
<intersection>-86.5 1</intersection>
<intersection>-77 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>230,-77,234.5,-77</points>
<connection>
<GID>195</GID>
<name>count_enable</name></connection>
<intersection>230 4</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>233.5,-86.5,233.5,-86</points>
<connection>
<GID>195</GID>
<name>clock</name></connection>
<intersection>-86.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,-43,302.5,-26</points>
<connection>
<GID>206</GID>
<name>IN_3</name></connection>
<intersection>-39 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>297,-39,302.5,-39</points>
<intersection>297 17</intersection>
<intersection>302.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301,-26,302.5,-26</points>
<connection>
<GID>207</GID>
<name>OUT_3</name></connection>
<intersection>302.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>297,-39,297,-38.5</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301,-46,301,-29</points>
<connection>
<GID>207</GID>
<name>OUT_0</name></connection>
<intersection>-46 5</intersection>
<intersection>-38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>299,-38.5,301,-38.5</points>
<connection>
<GID>208</GID>
<name>IN_1</name></connection>
<intersection>301 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>301,-46,302.5,-46</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>301 0</intersection></hsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-44,302,-27</points>
<intersection>-44 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302,-44,302.5,-44</points>
<connection>
<GID>206</GID>
<name>IN_2</name></connection>
<intersection>302 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301,-27,302,-27</points>
<connection>
<GID>207</GID>
<name>OUT_2</name></connection>
<intersection>302 0</intersection></hsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-45,301.5,-28</points>
<intersection>-45 3</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>301,-28,301.5,-28</points>
<connection>
<GID>207</GID>
<name>OUT_1</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>301.5,-45,302.5,-45</points>
<connection>
<GID>206</GID>
<name>IN_1</name></connection>
<intersection>301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298,-32.5,298,-32</points>
<connection>
<GID>208</GID>
<name>OUT</name></connection>
<connection>
<GID>207</GID>
<name>clear</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282,-32.5,298,-32.5</points>
<intersection>282 2</intersection>
<intersection>285.5 7</intersection>
<intersection>298 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>282,-32.5,282,-22.5</points>
<intersection>-32.5 1</intersection>
<intersection>-22.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>282,-22.5,286.5,-22.5</points>
<intersection>282 2</intersection>
<intersection>286.5 10</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>285.5,-32.5,285.5,-32</points>
<connection>
<GID>210</GID>
<name>clock</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>286.5,-23,286.5,-22.5</points>
<connection>
<GID>210</GID>
<name>count_enable</name></connection>
<intersection>-22.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,-43,292,-26</points>
<connection>
<GID>209</GID>
<name>IN_3</name></connection>
<intersection>-39 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286.5,-39,292,-39</points>
<intersection>286.5 17</intersection>
<intersection>292 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>290.5,-26,292,-26</points>
<connection>
<GID>210</GID>
<name>OUT_3</name></connection>
<intersection>292 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>286.5,-39,286.5,-38.5</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-46,290.5,-29</points>
<connection>
<GID>210</GID>
<name>OUT_0</name></connection>
<intersection>-46 5</intersection>
<intersection>-38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>288.5,-38.5,290.5,-38.5</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<intersection>290.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>290.5,-46,292,-46</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>290.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,-44,291.5,-27</points>
<intersection>-44 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>291.5,-44,292,-44</points>
<connection>
<GID>209</GID>
<name>IN_2</name></connection>
<intersection>291.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>290.5,-27,291.5,-27</points>
<connection>
<GID>210</GID>
<name>OUT_2</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,-45,291,-28</points>
<intersection>-45 3</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>290.5,-28,291,-28</points>
<connection>
<GID>210</GID>
<name>OUT_1</name></connection>
<intersection>291 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>291,-45,292,-45</points>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<intersection>291 0</intersection></hsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287.5,-32.5,287.5,-32</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<connection>
<GID>210</GID>
<name>clear</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>271.5,-32.5,287.5,-32.5</points>
<intersection>271.5 2</intersection>
<intersection>275 12</intersection>
<intersection>287.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>271.5,-32.5,271.5,-23</points>
<intersection>-32.5 1</intersection>
<intersection>-23 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>271.5,-23,276,-23</points>
<connection>
<GID>213</GID>
<name>count_enable</name></connection>
<intersection>271.5 2</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>275,-32.5,275,-32</points>
<connection>
<GID>213</GID>
<name>clock</name></connection>
<intersection>-32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-43,281.5,-26</points>
<connection>
<GID>212</GID>
<name>IN_3</name></connection>
<intersection>-39 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-39,281.5,-39</points>
<intersection>276 17</intersection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280,-26,281.5,-26</points>
<connection>
<GID>213</GID>
<name>OUT_3</name></connection>
<intersection>281.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>276,-39,276,-38.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280,-46,280,-29</points>
<connection>
<GID>213</GID>
<name>OUT_0</name></connection>
<intersection>-46 5</intersection>
<intersection>-38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>278,-38.5,280,-38.5</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<intersection>280 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>280,-46,281.5,-46</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>280 0</intersection></hsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,-44,281,-27</points>
<intersection>-44 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281,-44,281.5,-44</points>
<connection>
<GID>212</GID>
<name>IN_2</name></connection>
<intersection>281 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280,-27,281,-27</points>
<connection>
<GID>213</GID>
<name>OUT_2</name></connection>
<intersection>281 0</intersection></hsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280.5,-45,280.5,-28</points>
<intersection>-45 3</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>280,-28,280.5,-28</points>
<connection>
<GID>213</GID>
<name>OUT_1</name></connection>
<intersection>280.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>280.5,-45,281.5,-45</points>
<connection>
<GID>212</GID>
<name>IN_1</name></connection>
<intersection>280.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-43,271,-26</points>
<connection>
<GID>215</GID>
<name>IN_3</name></connection>
<intersection>-39 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>265.5,-39,271,-39</points>
<intersection>265.5 17</intersection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>269.5,-26,271,-26</points>
<connection>
<GID>246</GID>
<name>OUT_3</name></connection>
<intersection>271 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>265.5,-39,265.5,-38.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269.5,-46,269.5,-29</points>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection>
<intersection>-46 5</intersection>
<intersection>-38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>267.5,-38.5,269.5,-38.5</points>
<connection>
<GID>247</GID>
<name>IN_1</name></connection>
<intersection>269.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>269.5,-46,271,-46</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>269.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-44,270.5,-27</points>
<intersection>-44 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270.5,-44,271,-44</points>
<connection>
<GID>215</GID>
<name>IN_2</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>269.5,-27,270.5,-27</points>
<connection>
<GID>246</GID>
<name>OUT_2</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,-45,270,-28</points>
<intersection>-45 3</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>269.5,-28,270,-28</points>
<connection>
<GID>246</GID>
<name>OUT_1</name></connection>
<intersection>270 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>270,-45,271,-45</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<intersection>270 0</intersection></hsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,-32.5,261,-22.5</points>
<intersection>-32.5 4</intersection>
<intersection>-22.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>261,-22.5,265.5,-22.5</points>
<intersection>261 0</intersection>
<intersection>265.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>261,-32.5,277,-32.5</points>
<intersection>261 0</intersection>
<intersection>264.5 7</intersection>
<intersection>277 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>277,-32.5,277,-32</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<connection>
<GID>213</GID>
<name>clear</name></connection>
<intersection>-32.5 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>264.5,-32.5,264.5,-32</points>
<connection>
<GID>246</GID>
<name>clock</name></connection>
<intersection>-32.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>265.5,-23,265.5,-22.5</points>
<connection>
<GID>246</GID>
<name>count_enable</name></connection>
<intersection>-22.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,-43,260.5,-26</points>
<connection>
<GID>248</GID>
<name>IN_3</name></connection>
<intersection>-39 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255,-39,260.5,-39</points>
<intersection>255 17</intersection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259,-26,260.5,-26</points>
<connection>
<GID>249</GID>
<name>OUT_3</name></connection>
<intersection>260.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>255,-39,255,-38.5</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259,-46,259,-29</points>
<connection>
<GID>249</GID>
<name>OUT_0</name></connection>
<intersection>-46 5</intersection>
<intersection>-38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>257,-38.5,259,-38.5</points>
<connection>
<GID>250</GID>
<name>IN_1</name></connection>
<intersection>259 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>259,-46,260.5,-46</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>259 0</intersection></hsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-44,260,-27</points>
<intersection>-44 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,-44,260.5,-44</points>
<connection>
<GID>248</GID>
<name>IN_2</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259,-27,260,-27</points>
<connection>
<GID>249</GID>
<name>OUT_2</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,-45,259.5,-28</points>
<intersection>-45 3</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>259,-28,259.5,-28</points>
<connection>
<GID>249</GID>
<name>OUT_1</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>259.5,-45,260.5,-45</points>
<connection>
<GID>248</GID>
<name>IN_1</name></connection>
<intersection>259.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,-32,250.5,-22.5</points>
<intersection>-32 4</intersection>
<intersection>-22.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>250.5,-22.5,255,-22.5</points>
<intersection>250.5 0</intersection>
<intersection>255 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>250.5,-32,266.5,-32</points>
<connection>
<GID>249</GID>
<name>clock</name></connection>
<intersection>250.5 0</intersection>
<intersection>266.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>266.5,-32.5,266.5,-32</points>
<connection>
<GID>247</GID>
<name>OUT</name></connection>
<connection>
<GID>246</GID>
<name>clear</name></connection>
<intersection>-32 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>255,-23,255,-22.5</points>
<connection>
<GID>249</GID>
<name>count_enable</name></connection>
<intersection>-22.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,-32,292.5,-22</points>
<intersection>-32 4</intersection>
<intersection>-22 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>197,-22,297,-22</points>
<intersection>197 7</intersection>
<intersection>292.5 0</intersection>
<intersection>297 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>292.5,-32,296,-32</points>
<connection>
<GID>207</GID>
<name>clock</name></connection>
<intersection>292.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>297,-23,297,-22</points>
<connection>
<GID>207</GID>
<name>count_enable</name></connection>
<intersection>-22 3</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>197,-59.5,197,-22</points>
<intersection>-59.5 8</intersection>
<intersection>-22 3</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>197,-59.5,204,-59.5</points>
<connection>
<GID>184</GID>
<name>clear</name></connection>
<intersection>197 7</intersection>
<intersection>204 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>204,-60,204,-59.5</points>
<connection>
<GID>185</GID>
<name>OUT</name></connection>
<intersection>-59.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,-43,250,-26</points>
<connection>
<GID>251</GID>
<name>IN_3</name></connection>
<intersection>-39 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244.5,-39,250,-39</points>
<intersection>244.5 17</intersection>
<intersection>250 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>248.5,-26,250,-26</points>
<connection>
<GID>252</GID>
<name>OUT_3</name></connection>
<intersection>250 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>244.5,-39,244.5,-38.5</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,-16.5,302.5,0.5</points>
<connection>
<GID>216</GID>
<name>IN_3</name></connection>
<intersection>-12.5 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>297,-12.5,302.5,-12.5</points>
<intersection>297 17</intersection>
<intersection>302.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301,0.5,302.5,0.5</points>
<connection>
<GID>217</GID>
<name>OUT_3</name></connection>
<intersection>302.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>297,-12.5,297,-12</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>-12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301,-19.5,301,-2.5</points>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 5</intersection>
<intersection>-12 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>299,-12,301,-12</points>
<connection>
<GID>218</GID>
<name>IN_1</name></connection>
<intersection>301 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>301,-19.5,302.5,-19.5</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>301 0</intersection></hsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-17.5,302,-0.5</points>
<intersection>-17.5 1</intersection>
<intersection>-0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302,-17.5,302.5,-17.5</points>
<connection>
<GID>216</GID>
<name>IN_2</name></connection>
<intersection>302 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301,-0.5,302,-0.5</points>
<connection>
<GID>217</GID>
<name>OUT_2</name></connection>
<intersection>302 0</intersection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-18.5,301.5,-1.5</points>
<intersection>-18.5 3</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>301,-1.5,301.5,-1.5</points>
<connection>
<GID>217</GID>
<name>OUT_1</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>301.5,-18.5,302.5,-18.5</points>
<connection>
<GID>216</GID>
<name>IN_1</name></connection>
<intersection>301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298,-6,298,-5.5</points>
<connection>
<GID>218</GID>
<name>OUT</name></connection>
<connection>
<GID>217</GID>
<name>clear</name></connection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282,-6,298,-6</points>
<intersection>282 2</intersection>
<intersection>285.5 7</intersection>
<intersection>298 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>282,-6,282,4</points>
<intersection>-6 1</intersection>
<intersection>4 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>282,4,286.5,4</points>
<intersection>282 2</intersection>
<intersection>286.5 10</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>285.5,-6,285.5,-5.5</points>
<connection>
<GID>220</GID>
<name>clock</name></connection>
<intersection>-6 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>286.5,3.5,286.5,4</points>
<connection>
<GID>220</GID>
<name>count_enable</name></connection>
<intersection>4 5</intersection></vsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248.5,-46,248.5,-29</points>
<connection>
<GID>252</GID>
<name>OUT_0</name></connection>
<intersection>-46 5</intersection>
<intersection>-38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>246.5,-38.5,248.5,-38.5</points>
<connection>
<GID>253</GID>
<name>IN_1</name></connection>
<intersection>248.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>248.5,-46,250,-46</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>248.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,-16.5,292,0.5</points>
<connection>
<GID>219</GID>
<name>IN_3</name></connection>
<intersection>-12.5 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286.5,-12.5,292,-12.5</points>
<intersection>286.5 17</intersection>
<intersection>292 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>290.5,0.5,292,0.5</points>
<connection>
<GID>220</GID>
<name>OUT_3</name></connection>
<intersection>292 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>286.5,-12.5,286.5,-12</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>-12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-19.5,290.5,-2.5</points>
<connection>
<GID>220</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 5</intersection>
<intersection>-12 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>288.5,-12,290.5,-12</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<intersection>290.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>290.5,-19.5,292,-19.5</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>290.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,-17.5,291.5,-0.5</points>
<intersection>-17.5 1</intersection>
<intersection>-0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>291.5,-17.5,292,-17.5</points>
<connection>
<GID>219</GID>
<name>IN_2</name></connection>
<intersection>291.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>290.5,-0.5,291.5,-0.5</points>
<connection>
<GID>220</GID>
<name>OUT_2</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,-18.5,291,-1.5</points>
<intersection>-18.5 3</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>290.5,-1.5,291,-1.5</points>
<connection>
<GID>220</GID>
<name>OUT_1</name></connection>
<intersection>291 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>291,-18.5,292,-18.5</points>
<connection>
<GID>219</GID>
<name>IN_1</name></connection>
<intersection>291 0</intersection></hsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287.5,-6,287.5,-5.5</points>
<connection>
<GID>221</GID>
<name>OUT</name></connection>
<connection>
<GID>220</GID>
<name>clear</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>271.5,-5.5,287.5,-5.5</points>
<connection>
<GID>223</GID>
<name>clock</name></connection>
<intersection>271.5 2</intersection>
<intersection>287.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>271.5,-5.5,271.5,4</points>
<intersection>-5.5 1</intersection>
<intersection>4 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>271.5,4,276,4</points>
<intersection>271.5 2</intersection>
<intersection>276 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>276,3.5,276,4</points>
<connection>
<GID>223</GID>
<name>count_enable</name></connection>
<intersection>4 5</intersection></vsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-16.5,281.5,0.5</points>
<connection>
<GID>222</GID>
<name>IN_3</name></connection>
<intersection>-12.5 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-12.5,281.5,-12.5</points>
<intersection>276 17</intersection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280,0.5,281.5,0.5</points>
<connection>
<GID>223</GID>
<name>OUT_3</name></connection>
<intersection>281.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>276,-12.5,276,-12</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>-12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280,-19.5,280,-2.5</points>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 5</intersection>
<intersection>-12 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>278,-12,280,-12</points>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<intersection>280 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>280,-19.5,281.5,-19.5</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>280 0</intersection></hsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,-17.5,281,-0.5</points>
<intersection>-17.5 1</intersection>
<intersection>-0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281,-17.5,281.5,-17.5</points>
<connection>
<GID>222</GID>
<name>IN_2</name></connection>
<intersection>281 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280,-0.5,281,-0.5</points>
<connection>
<GID>223</GID>
<name>OUT_2</name></connection>
<intersection>281 0</intersection></hsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280.5,-18.5,280.5,-1.5</points>
<intersection>-18.5 3</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>280,-1.5,280.5,-1.5</points>
<connection>
<GID>223</GID>
<name>OUT_1</name></connection>
<intersection>280.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>280.5,-18.5,281.5,-18.5</points>
<connection>
<GID>222</GID>
<name>IN_1</name></connection>
<intersection>280.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-16.5,271,0.5</points>
<connection>
<GID>225</GID>
<name>IN_3</name></connection>
<intersection>-12.5 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>265.5,-12.5,271,-12.5</points>
<intersection>265.5 17</intersection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>269.5,0.5,271,0.5</points>
<connection>
<GID>226</GID>
<name>OUT_3</name></connection>
<intersection>271 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>265.5,-12.5,265.5,-12</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>-12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269.5,-19.5,269.5,-2.5</points>
<connection>
<GID>226</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 5</intersection>
<intersection>-12 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>267.5,-12,269.5,-12</points>
<connection>
<GID>227</GID>
<name>IN_1</name></connection>
<intersection>269.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>269.5,-19.5,271,-19.5</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>269.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-17.5,270.5,-0.5</points>
<intersection>-17.5 1</intersection>
<intersection>-0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270.5,-17.5,271,-17.5</points>
<connection>
<GID>225</GID>
<name>IN_2</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>269.5,-0.5,270.5,-0.5</points>
<connection>
<GID>226</GID>
<name>OUT_2</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,-18.5,270,-1.5</points>
<intersection>-18.5 3</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>269.5,-1.5,270,-1.5</points>
<connection>
<GID>226</GID>
<name>OUT_1</name></connection>
<intersection>270 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>270,-18.5,271,-18.5</points>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<intersection>270 0</intersection></hsegment></shape></wire>
<wire>
<ID>386</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,-6,261,4</points>
<intersection>-6 4</intersection>
<intersection>4 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>261,4,265.5,4</points>
<intersection>261 0</intersection>
<intersection>265.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>261,-6,277,-6</points>
<intersection>261 0</intersection>
<intersection>264.5 7</intersection>
<intersection>277 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>277,-6,277,-5.5</points>
<connection>
<GID>224</GID>
<name>OUT</name></connection>
<connection>
<GID>223</GID>
<name>clear</name></connection>
<intersection>-6 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>264.5,-6,264.5,-5.5</points>
<connection>
<GID>226</GID>
<name>clock</name></connection>
<intersection>-6 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>265.5,3.5,265.5,4</points>
<connection>
<GID>226</GID>
<name>count_enable</name></connection>
<intersection>4 3</intersection></vsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,-16.5,260.5,0.5</points>
<connection>
<GID>228</GID>
<name>IN_3</name></connection>
<intersection>-12.5 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255,-12.5,260.5,-12.5</points>
<intersection>255 17</intersection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259,0.5,260.5,0.5</points>
<connection>
<GID>229</GID>
<name>OUT_3</name></connection>
<intersection>260.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>255,-12.5,255,-12</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>-12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259,-19.5,259,-2.5</points>
<connection>
<GID>229</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 5</intersection>
<intersection>-12 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>257,-12,259,-12</points>
<connection>
<GID>230</GID>
<name>IN_1</name></connection>
<intersection>259 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>259,-19.5,260.5,-19.5</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>259 0</intersection></hsegment></shape></wire>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-17.5,260,-0.5</points>
<intersection>-17.5 1</intersection>
<intersection>-0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,-17.5,260.5,-17.5</points>
<connection>
<GID>228</GID>
<name>IN_2</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259,-0.5,260,-0.5</points>
<connection>
<GID>229</GID>
<name>OUT_2</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,-18.5,259.5,-1.5</points>
<intersection>-18.5 3</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>259,-1.5,259.5,-1.5</points>
<connection>
<GID>229</GID>
<name>OUT_1</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>259.5,-18.5,260.5,-18.5</points>
<connection>
<GID>228</GID>
<name>IN_1</name></connection>
<intersection>259.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,-44,249.5,-27</points>
<intersection>-44 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>249.5,-44,250,-44</points>
<connection>
<GID>251</GID>
<name>IN_2</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>248.5,-27,249.5,-27</points>
<connection>
<GID>252</GID>
<name>OUT_2</name></connection>
<intersection>249.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,-5.5,250.5,4</points>
<intersection>-5.5 4</intersection>
<intersection>4 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>250.5,4,255,4</points>
<intersection>250.5 0</intersection>
<intersection>255 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>250.5,-5.5,266.5,-5.5</points>
<connection>
<GID>229</GID>
<name>clock</name></connection>
<intersection>250.5 0</intersection>
<intersection>266.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>266.5,-6,266.5,-5.5</points>
<connection>
<GID>227</GID>
<name>OUT</name></connection>
<connection>
<GID>226</GID>
<name>clear</name></connection>
<intersection>-5.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>255,3.5,255,4</points>
<connection>
<GID>229</GID>
<name>count_enable</name></connection>
<intersection>4 3</intersection></vsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,-5.5,292.5,4</points>
<intersection>-5.5 4</intersection>
<intersection>4 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>292.5,4,297,4</points>
<intersection>292.5 0</intersection>
<intersection>297 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>292.5,-5.5,296,-5.5</points>
<connection>
<GID>217</GID>
<name>clock</name></connection>
<intersection>292.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>297,3.5,297,5</points>
<connection>
<GID>217</GID>
<name>count_enable</name></connection>
<intersection>4 3</intersection>
<intersection>5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>196,5,297,5</points>
<intersection>196 7</intersection>
<intersection>297 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>196,-32.5,196,5</points>
<intersection>-32.5 8</intersection>
<intersection>5 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>196,-32.5,203.5,-32.5</points>
<connection>
<GID>265</GID>
<name>OUT</name></connection>
<intersection>196 7</intersection>
<intersection>203.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>203.5,-32.5,203.5,-32</points>
<connection>
<GID>264</GID>
<name>clear</name></connection>
<intersection>-32.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,-16.5,250,0.5</points>
<connection>
<GID>231</GID>
<name>IN_3</name></connection>
<intersection>-12.5 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244.5,-12.5,250,-12.5</points>
<intersection>244.5 17</intersection>
<intersection>250 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>248.5,0.5,250,0.5</points>
<connection>
<GID>232</GID>
<name>OUT_3</name></connection>
<intersection>250 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>244.5,-12.5,244.5,-12</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>-12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248.5,-19.5,248.5,-2.5</points>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 5</intersection>
<intersection>-12 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>246.5,-12,248.5,-12</points>
<connection>
<GID>233</GID>
<name>IN_1</name></connection>
<intersection>248.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>248.5,-19.5,250,-19.5</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>248.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,-17.5,249.5,-0.5</points>
<intersection>-17.5 1</intersection>
<intersection>-0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>249.5,-17.5,250,-17.5</points>
<connection>
<GID>231</GID>
<name>IN_2</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>248.5,-0.5,249.5,-0.5</points>
<connection>
<GID>232</GID>
<name>OUT_2</name></connection>
<intersection>249.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249,-18.5,249,-1.5</points>
<intersection>-18.5 3</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>248.5,-1.5,249,-1.5</points>
<connection>
<GID>232</GID>
<name>OUT_1</name></connection>
<intersection>249 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>249,-18.5,250,-18.5</points>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<intersection>249 0</intersection></hsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249,-45,249,-28</points>
<intersection>-45 3</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>248.5,-28,249,-28</points>
<connection>
<GID>252</GID>
<name>OUT_1</name></connection>
<intersection>249 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>249,-45,250,-45</points>
<connection>
<GID>251</GID>
<name>IN_1</name></connection>
<intersection>249 0</intersection></hsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239.5,-16.5,239.5,0.5</points>
<connection>
<GID>234</GID>
<name>IN_3</name></connection>
<intersection>-12.5 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234,-12.5,239.5,-12.5</points>
<intersection>234 17</intersection>
<intersection>239.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238,0.5,239.5,0.5</points>
<connection>
<GID>235</GID>
<name>OUT_3</name></connection>
<intersection>239.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>234,-12.5,234,-12</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>-12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238,-19.5,238,-2.5</points>
<connection>
<GID>235</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 5</intersection>
<intersection>-12 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>236,-12,238,-12</points>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>238,-19.5,239.5,-19.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>238 0</intersection></hsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,-17.5,239,-0.5</points>
<intersection>-17.5 1</intersection>
<intersection>-0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239,-17.5,239.5,-17.5</points>
<connection>
<GID>234</GID>
<name>IN_2</name></connection>
<intersection>239 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238,-0.5,239,-0.5</points>
<connection>
<GID>235</GID>
<name>OUT_2</name></connection>
<intersection>239 0</intersection></hsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,-18.5,238.5,-1.5</points>
<intersection>-18.5 3</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>238,-1.5,238.5,-1.5</points>
<connection>
<GID>235</GID>
<name>OUT_1</name></connection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>238.5,-18.5,239.5,-18.5</points>
<connection>
<GID>234</GID>
<name>IN_1</name></connection>
<intersection>238.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,-6,235,-5.5</points>
<connection>
<GID>236</GID>
<name>OUT</name></connection>
<connection>
<GID>235</GID>
<name>clear</name></connection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,-6,235,-6</points>
<intersection>219 2</intersection>
<intersection>222.5 10</intersection>
<intersection>235 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>219,-6,219,4</points>
<intersection>-6 1</intersection>
<intersection>4 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>219,4,223.5,4</points>
<intersection>219 2</intersection>
<intersection>223.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>223.5,3.5,223.5,4</points>
<connection>
<GID>238</GID>
<name>count_enable</name></connection>
<intersection>4 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>222.5,-6,222.5,-5.5</points>
<connection>
<GID>238</GID>
<name>clock</name></connection>
<intersection>-6 1</intersection></vsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-16.5,229,0.5</points>
<connection>
<GID>237</GID>
<name>IN_3</name></connection>
<intersection>-12.5 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>223.5,-12.5,229,-12.5</points>
<intersection>223.5 17</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227.5,0.5,229,0.5</points>
<connection>
<GID>238</GID>
<name>OUT_3</name></connection>
<intersection>229 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>223.5,-12.5,223.5,-12</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>-12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227.5,-19.5,227.5,-2.5</points>
<connection>
<GID>238</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 5</intersection>
<intersection>-12 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>225.5,-12,227.5,-12</points>
<connection>
<GID>239</GID>
<name>IN_1</name></connection>
<intersection>227.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>227.5,-19.5,229,-19.5</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>227.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,-17.5,228.5,-0.5</points>
<intersection>-17.5 1</intersection>
<intersection>-0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>228.5,-17.5,229,-17.5</points>
<connection>
<GID>237</GID>
<name>IN_2</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227.5,-0.5,228.5,-0.5</points>
<connection>
<GID>238</GID>
<name>OUT_2</name></connection>
<intersection>228.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,-18.5,228,-1.5</points>
<intersection>-18.5 3</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>227.5,-1.5,228,-1.5</points>
<connection>
<GID>238</GID>
<name>OUT_1</name></connection>
<intersection>228 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>228,-18.5,229,-18.5</points>
<connection>
<GID>237</GID>
<name>IN_1</name></connection>
<intersection>228 0</intersection></hsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-16.5,218.5,0.5</points>
<connection>
<GID>240</GID>
<name>IN_3</name></connection>
<intersection>-12.5 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213,-12.5,218.5,-12.5</points>
<intersection>213 17</intersection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>217,0.5,218.5,0.5</points>
<connection>
<GID>241</GID>
<name>OUT_3</name></connection>
<intersection>218.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>213,-12.5,213,-12</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>-12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217,-19.5,217,-2.5</points>
<connection>
<GID>241</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 5</intersection>
<intersection>-12 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>215,-12,217,-12</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>217,-19.5,218.5,-19.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-17.5,218,-0.5</points>
<intersection>-17.5 1</intersection>
<intersection>-0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,-17.5,218.5,-17.5</points>
<connection>
<GID>240</GID>
<name>IN_2</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>217,-0.5,218,-0.5</points>
<connection>
<GID>241</GID>
<name>OUT_2</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217.5,-18.5,217.5,-1.5</points>
<intersection>-18.5 3</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>217,-1.5,217.5,-1.5</points>
<connection>
<GID>241</GID>
<name>OUT_1</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>217.5,-18.5,218.5,-18.5</points>
<connection>
<GID>240</GID>
<name>IN_1</name></connection>
<intersection>217.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-5.5,208.5,4</points>
<intersection>-5.5 4</intersection>
<intersection>4 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>208.5,4,213,4</points>
<intersection>208.5 0</intersection>
<intersection>213 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>208.5,-5.5,224.5,-5.5</points>
<connection>
<GID>241</GID>
<name>clock</name></connection>
<intersection>208.5 0</intersection>
<intersection>224.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>224.5,-6,224.5,-5.5</points>
<connection>
<GID>239</GID>
<name>OUT</name></connection>
<connection>
<GID>238</GID>
<name>clear</name></connection>
<intersection>-5.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>213,3.5,213,4</points>
<connection>
<GID>241</GID>
<name>count_enable</name></connection>
<intersection>4 3</intersection></vsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-16.5,208,0.5</points>
<connection>
<GID>243</GID>
<name>IN_3</name></connection>
<intersection>-12.5 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,-12.5,208,-12.5</points>
<intersection>202.5 17</intersection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>206.5,0.5,208,0.5</points>
<connection>
<GID>244</GID>
<name>OUT_3</name></connection>
<intersection>208 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>202.5,-12.5,202.5,-12</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<intersection>-12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,-19.5,206.5,-2.5</points>
<connection>
<GID>244</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 5</intersection>
<intersection>-12 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>204.5,-12,206.5,-12</points>
<connection>
<GID>245</GID>
<name>IN_1</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>206.5,-19.5,208,-19.5</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>206.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,-17.5,207.5,-0.5</points>
<intersection>-17.5 1</intersection>
<intersection>-0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207.5,-17.5,208,-17.5</points>
<connection>
<GID>243</GID>
<name>IN_2</name></connection>
<intersection>207.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>206.5,-0.5,207.5,-0.5</points>
<connection>
<GID>244</GID>
<name>OUT_2</name></connection>
<intersection>207.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-18.5,207,-1.5</points>
<intersection>-18.5 3</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>206.5,-1.5,207,-1.5</points>
<connection>
<GID>244</GID>
<name>OUT_1</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>207,-18.5,208,-18.5</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203.5,-6,203.5,-5.5</points>
<connection>
<GID>245</GID>
<name>OUT</name></connection>
<connection>
<GID>244</GID>
<name>clear</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>197,-5.5,203.5,-5.5</points>
<intersection>197 2</intersection>
<intersection>203.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-5.5,197,31.5</points>
<intersection>-5.5 1</intersection>
<intersection>31.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>197,31.5,297,31.5</points>
<intersection>197 2</intersection>
<intersection>296 8</intersection>
<intersection>297 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>297,30.5,297,31.5</points>
<connection>
<GID>267</GID>
<name>count_enable</name></connection>
<intersection>31.5 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>296,21.5,296,31.5</points>
<connection>
<GID>267</GID>
<name>clock</name></connection>
<intersection>31.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198,-6,198,4</points>
<intersection>-6 4</intersection>
<intersection>4 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,4,202.5,4</points>
<intersection>198 0</intersection>
<intersection>202.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>198,-6,214,-6</points>
<intersection>198 0</intersection>
<intersection>201.5 15</intersection>
<intersection>214 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>214,-6,214,-5.5</points>
<connection>
<GID>242</GID>
<name>OUT</name></connection>
<connection>
<GID>241</GID>
<name>clear</name></connection>
<intersection>-6 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>202.5,3.5,202.5,4</points>
<connection>
<GID>244</GID>
<name>count_enable</name></connection>
<intersection>4 3</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>201.5,-6,201.5,-5.5</points>
<connection>
<GID>244</GID>
<name>clock</name></connection>
<intersection>-6 4</intersection></vsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239.5,-43,239.5,-26</points>
<connection>
<GID>254</GID>
<name>IN_3</name></connection>
<intersection>-39 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234,-39,239.5,-39</points>
<intersection>234 17</intersection>
<intersection>239.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238,-26,239.5,-26</points>
<connection>
<GID>255</GID>
<name>OUT_3</name></connection>
<intersection>239.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>234,-39,234,-38.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>256,-6,256,-5.5</points>
<connection>
<GID>230</GID>
<name>OUT</name></connection>
<connection>
<GID>229</GID>
<name>clear</name></connection>
<intersection>-6 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>240,-6,256,-6</points>
<intersection>240 4</intersection>
<intersection>243.5 8</intersection>
<intersection>256 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>240,-6,240,4</points>
<intersection>-6 3</intersection>
<intersection>4 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>240,4,244.5,4</points>
<intersection>240 4</intersection>
<intersection>244.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>244.5,3.5,244.5,4</points>
<connection>
<GID>232</GID>
<name>count_enable</name></connection>
<intersection>4 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>243.5,-6,243.5,-5.5</points>
<connection>
<GID>232</GID>
<name>clock</name></connection>
<intersection>-6 3</intersection></vsegment></shape></wire>
<wire>
<ID>421</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-6,245.5,-5.5</points>
<connection>
<GID>233</GID>
<name>OUT</name></connection>
<connection>
<GID>232</GID>
<name>clear</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229.5,-5.5,245.5,-5.5</points>
<connection>
<GID>235</GID>
<name>clock</name></connection>
<intersection>229.5 4</intersection>
<intersection>245.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>229.5,-5.5,229.5,4</points>
<intersection>-5.5 1</intersection>
<intersection>4 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>229.5,4,234,4</points>
<intersection>229.5 4</intersection>
<intersection>234 17</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>234,3.5,234,4</points>
<connection>
<GID>235</GID>
<name>count_enable</name></connection>
<intersection>4 15</intersection></vsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238,-46,238,-29</points>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection>
<intersection>-46 5</intersection>
<intersection>-38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>236,-38.5,238,-38.5</points>
<connection>
<GID>256</GID>
<name>IN_1</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>238,-46,239.5,-46</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>238 0</intersection></hsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,-44,239,-27</points>
<intersection>-44 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239,-44,239.5,-44</points>
<connection>
<GID>254</GID>
<name>IN_2</name></connection>
<intersection>239 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238,-27,239,-27</points>
<connection>
<GID>255</GID>
<name>OUT_2</name></connection>
<intersection>239 0</intersection></hsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,-45,238.5,-28</points>
<intersection>-45 3</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>238,-28,238.5,-28</points>
<connection>
<GID>255</GID>
<name>OUT_1</name></connection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>238.5,-45,239.5,-45</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<intersection>238.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,-32.5,235,-32</points>
<connection>
<GID>256</GID>
<name>OUT</name></connection>
<connection>
<GID>255</GID>
<name>clear</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,-32.5,235,-32.5</points>
<intersection>219 2</intersection>
<intersection>222.5 10</intersection>
<intersection>235 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>219,-32.5,219,-22.5</points>
<intersection>-32.5 1</intersection>
<intersection>-22.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>219,-22.5,223.5,-22.5</points>
<intersection>219 2</intersection>
<intersection>223.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>223.5,-23,223.5,-22.5</points>
<connection>
<GID>258</GID>
<name>count_enable</name></connection>
<intersection>-22.5 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>222.5,-32.5,222.5,-32</points>
<connection>
<GID>258</GID>
<name>clock</name></connection>
<intersection>-32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-43,229,-26</points>
<connection>
<GID>257</GID>
<name>IN_3</name></connection>
<intersection>-39 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>223.5,-39,229,-39</points>
<intersection>223.5 17</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227.5,-26,229,-26</points>
<connection>
<GID>258</GID>
<name>OUT_3</name></connection>
<intersection>229 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>223.5,-39,223.5,-38.5</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227.5,-46,227.5,-29</points>
<connection>
<GID>258</GID>
<name>OUT_0</name></connection>
<intersection>-46 5</intersection>
<intersection>-38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>225.5,-38.5,227.5,-38.5</points>
<connection>
<GID>259</GID>
<name>IN_1</name></connection>
<intersection>227.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>227.5,-46,229,-46</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>227.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,-44,228.5,-27</points>
<intersection>-44 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>228.5,-44,229,-44</points>
<connection>
<GID>257</GID>
<name>IN_2</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227.5,-27,228.5,-27</points>
<connection>
<GID>258</GID>
<name>OUT_2</name></connection>
<intersection>228.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,-45,228,-28</points>
<intersection>-45 3</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>227.5,-28,228,-28</points>
<connection>
<GID>258</GID>
<name>OUT_1</name></connection>
<intersection>228 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>228,-45,229,-45</points>
<connection>
<GID>257</GID>
<name>IN_1</name></connection>
<intersection>228 0</intersection></hsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-43,218.5,-26</points>
<connection>
<GID>260</GID>
<name>IN_3</name></connection>
<intersection>-39 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213,-39,218.5,-39</points>
<intersection>213 17</intersection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>217,-26,218.5,-26</points>
<connection>
<GID>261</GID>
<name>OUT_3</name></connection>
<intersection>218.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>213,-39,213,-38.5</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217,-46,217,-29</points>
<connection>
<GID>261</GID>
<name>OUT_0</name></connection>
<intersection>-46 5</intersection>
<intersection>-38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>215,-38.5,217,-38.5</points>
<connection>
<GID>262</GID>
<name>IN_1</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>217,-46,218.5,-46</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-44,218,-27</points>
<intersection>-44 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,-44,218.5,-44</points>
<connection>
<GID>260</GID>
<name>IN_2</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>217,-27,218,-27</points>
<connection>
<GID>261</GID>
<name>OUT_2</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217.5,-45,217.5,-28</points>
<intersection>-45 3</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>217,-28,217.5,-28</points>
<connection>
<GID>261</GID>
<name>OUT_1</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>217.5,-45,218.5,-45</points>
<connection>
<GID>260</GID>
<name>IN_1</name></connection>
<intersection>217.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-32,208.5,-22.5</points>
<intersection>-32 4</intersection>
<intersection>-22.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>208.5,-22.5,213,-22.5</points>
<intersection>208.5 0</intersection>
<intersection>213 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>208.5,-32,224.5,-32</points>
<connection>
<GID>261</GID>
<name>clock</name></connection>
<intersection>208.5 0</intersection>
<intersection>224.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>224.5,-32.5,224.5,-32</points>
<connection>
<GID>259</GID>
<name>OUT</name></connection>
<connection>
<GID>258</GID>
<name>clear</name></connection>
<intersection>-32 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>213,-23,213,-22.5</points>
<connection>
<GID>261</GID>
<name>count_enable</name></connection>
<intersection>-22.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-43,208,-26</points>
<connection>
<GID>263</GID>
<name>IN_3</name></connection>
<intersection>-39 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,-39,208,-39</points>
<intersection>202.5 17</intersection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>206.5,-26,208,-26</points>
<connection>
<GID>264</GID>
<name>OUT_3</name></connection>
<intersection>208 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>202.5,-39,202.5,-38.5</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,-46,206.5,-29</points>
<connection>
<GID>264</GID>
<name>OUT_0</name></connection>
<intersection>-46 5</intersection>
<intersection>-38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>204.5,-38.5,206.5,-38.5</points>
<connection>
<GID>265</GID>
<name>IN_1</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>206.5,-46,208,-46</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>206.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,-44,207.5,-27</points>
<intersection>-44 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207.5,-44,208,-44</points>
<connection>
<GID>263</GID>
<name>IN_2</name></connection>
<intersection>207.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>206.5,-27,207.5,-27</points>
<connection>
<GID>264</GID>
<name>OUT_2</name></connection>
<intersection>207.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-45,207,-28</points>
<intersection>-45 3</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>206.5,-28,207,-28</points>
<connection>
<GID>264</GID>
<name>OUT_1</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>207,-45,208,-45</points>
<connection>
<GID>263</GID>
<name>IN_1</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>439</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198,-32.5,198,-22.5</points>
<intersection>-32.5 4</intersection>
<intersection>-22.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-22.5,202.5,-22.5</points>
<intersection>198 0</intersection>
<intersection>202.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>198,-32.5,214,-32.5</points>
<intersection>198 0</intersection>
<intersection>201.5 15</intersection>
<intersection>214 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>214,-32.5,214,-32</points>
<connection>
<GID>262</GID>
<name>OUT</name></connection>
<connection>
<GID>261</GID>
<name>clear</name></connection>
<intersection>-32.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>202.5,-23,202.5,-22.5</points>
<connection>
<GID>264</GID>
<name>count_enable</name></connection>
<intersection>-22.5 3</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>201.5,-32.5,201.5,-32</points>
<connection>
<GID>264</GID>
<name>clock</name></connection>
<intersection>-32.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>256,-32.5,256,-32</points>
<connection>
<GID>250</GID>
<name>OUT</name></connection>
<connection>
<GID>249</GID>
<name>clear</name></connection>
<intersection>-32.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>240,-32.5,256,-32.5</points>
<intersection>240 4</intersection>
<intersection>243.5 8</intersection>
<intersection>256 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>240,-32.5,240,-22.5</points>
<intersection>-32.5 3</intersection>
<intersection>-22.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>240,-22.5,244.5,-22.5</points>
<intersection>240 4</intersection>
<intersection>244.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>244.5,-23,244.5,-22.5</points>
<connection>
<GID>252</GID>
<name>count_enable</name></connection>
<intersection>-22.5 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>243.5,-32.5,243.5,-32</points>
<connection>
<GID>252</GID>
<name>clock</name></connection>
<intersection>-32.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>441</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-32.5,245.5,-32</points>
<connection>
<GID>253</GID>
<name>OUT</name></connection>
<connection>
<GID>252</GID>
<name>clear</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229.5,-32.5,245.5,-32.5</points>
<intersection>229.5 4</intersection>
<intersection>233 20</intersection>
<intersection>245.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>229.5,-32.5,229.5,-23</points>
<intersection>-32.5 1</intersection>
<intersection>-23 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>229.5,-23,234,-23</points>
<connection>
<GID>255</GID>
<name>count_enable</name></connection>
<intersection>229.5 4</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>233,-32.5,233,-32</points>
<connection>
<GID>255</GID>
<name>clock</name></connection>
<intersection>-32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,10.5,302.5,27.5</points>
<connection>
<GID>266</GID>
<name>IN_3</name></connection>
<intersection>14.5 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>297,14.5,302.5,14.5</points>
<intersection>297 17</intersection>
<intersection>302.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301,27.5,302.5,27.5</points>
<connection>
<GID>267</GID>
<name>OUT_3</name></connection>
<intersection>302.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>297,14.5,297,15</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>443</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301,7.5,301,24.5</points>
<connection>
<GID>267</GID>
<name>OUT_0</name></connection>
<intersection>7.5 5</intersection>
<intersection>15 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>299,15,301,15</points>
<connection>
<GID>268</GID>
<name>IN_1</name></connection>
<intersection>301 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>301,7.5,302.5,7.5</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>301 0</intersection></hsegment></shape></wire>
<wire>
<ID>444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,9.5,302,26.5</points>
<intersection>9.5 1</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302,9.5,302.5,9.5</points>
<connection>
<GID>266</GID>
<name>IN_2</name></connection>
<intersection>302 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301,26.5,302,26.5</points>
<connection>
<GID>267</GID>
<name>OUT_2</name></connection>
<intersection>302 0</intersection></hsegment></shape></wire>
<wire>
<ID>445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,8.5,301.5,25.5</points>
<intersection>8.5 3</intersection>
<intersection>25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>301,25.5,301.5,25.5</points>
<connection>
<GID>267</GID>
<name>OUT_1</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>301.5,8.5,302.5,8.5</points>
<connection>
<GID>266</GID>
<name>IN_1</name></connection>
<intersection>301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>446</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298,21,298,21.5</points>
<connection>
<GID>268</GID>
<name>OUT</name></connection>
<connection>
<GID>267</GID>
<name>clear</name></connection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282,21,298,21</points>
<intersection>282 2</intersection>
<intersection>285.5 7</intersection>
<intersection>298 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>282,21,282,31</points>
<intersection>21 1</intersection>
<intersection>31 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>282,31,286.5,31</points>
<intersection>282 2</intersection>
<intersection>286.5 10</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>285.5,21,285.5,21.5</points>
<connection>
<GID>270</GID>
<name>clock</name></connection>
<intersection>21 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>286.5,30.5,286.5,31</points>
<connection>
<GID>270</GID>
<name>count_enable</name></connection>
<intersection>31 5</intersection></vsegment></shape></wire>
<wire>
<ID>447</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,10.5,292,27.5</points>
<connection>
<GID>269</GID>
<name>IN_3</name></connection>
<intersection>14.5 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286.5,14.5,292,14.5</points>
<intersection>286.5 17</intersection>
<intersection>292 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>290.5,27.5,292,27.5</points>
<connection>
<GID>270</GID>
<name>OUT_3</name></connection>
<intersection>292 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>286.5,14.5,286.5,15</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>448</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,7.5,290.5,24.5</points>
<connection>
<GID>270</GID>
<name>OUT_0</name></connection>
<intersection>7.5 5</intersection>
<intersection>15 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>288.5,15,290.5,15</points>
<connection>
<GID>271</GID>
<name>IN_1</name></connection>
<intersection>290.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>290.5,7.5,292,7.5</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>290.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>449</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,9.5,291.5,26.5</points>
<intersection>9.5 1</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>291.5,9.5,292,9.5</points>
<connection>
<GID>269</GID>
<name>IN_2</name></connection>
<intersection>291.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>290.5,26.5,291.5,26.5</points>
<connection>
<GID>270</GID>
<name>OUT_2</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>450</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,8.5,291,25.5</points>
<intersection>8.5 3</intersection>
<intersection>25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>290.5,25.5,291,25.5</points>
<connection>
<GID>270</GID>
<name>OUT_1</name></connection>
<intersection>291 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>291,8.5,292,8.5</points>
<connection>
<GID>269</GID>
<name>IN_1</name></connection>
<intersection>291 0</intersection></hsegment></shape></wire>
<wire>
<ID>451</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287.5,21,287.5,21.5</points>
<connection>
<GID>271</GID>
<name>OUT</name></connection>
<connection>
<GID>270</GID>
<name>clear</name></connection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>271.5,21,287.5,21</points>
<intersection>271.5 2</intersection>
<intersection>275 12</intersection>
<intersection>287.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>271.5,21,271.5,30.5</points>
<intersection>21 1</intersection>
<intersection>30.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>271.5,30.5,276,30.5</points>
<connection>
<GID>273</GID>
<name>count_enable</name></connection>
<intersection>271.5 2</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>275,21,275,21.5</points>
<connection>
<GID>273</GID>
<name>clock</name></connection>
<intersection>21 1</intersection></vsegment></shape></wire>
<wire>
<ID>452</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,10.5,281.5,27.5</points>
<connection>
<GID>272</GID>
<name>IN_3</name></connection>
<intersection>14.5 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,14.5,281.5,14.5</points>
<intersection>276 17</intersection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280,27.5,281.5,27.5</points>
<connection>
<GID>273</GID>
<name>OUT_3</name></connection>
<intersection>281.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>276,14.5,276,15</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>453</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280,7.5,280,24.5</points>
<connection>
<GID>273</GID>
<name>OUT_0</name></connection>
<intersection>7.5 5</intersection>
<intersection>15 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>278,15,280,15</points>
<connection>
<GID>274</GID>
<name>IN_1</name></connection>
<intersection>280 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>280,7.5,281.5,7.5</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>280 0</intersection></hsegment></shape></wire>
<wire>
<ID>454</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,9.5,281,26.5</points>
<intersection>9.5 1</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281,9.5,281.5,9.5</points>
<connection>
<GID>272</GID>
<name>IN_2</name></connection>
<intersection>281 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280,26.5,281,26.5</points>
<connection>
<GID>273</GID>
<name>OUT_2</name></connection>
<intersection>281 0</intersection></hsegment></shape></wire>
<wire>
<ID>455</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280.5,8.5,280.5,25.5</points>
<intersection>8.5 3</intersection>
<intersection>25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>280,25.5,280.5,25.5</points>
<connection>
<GID>273</GID>
<name>OUT_1</name></connection>
<intersection>280.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>280.5,8.5,281.5,8.5</points>
<connection>
<GID>272</GID>
<name>IN_1</name></connection>
<intersection>280.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,10.5,271,27.5</points>
<connection>
<GID>275</GID>
<name>IN_3</name></connection>
<intersection>14.5 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>265.5,14.5,271,14.5</points>
<intersection>265.5 17</intersection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>269.5,27.5,271,27.5</points>
<connection>
<GID>306</GID>
<name>OUT_3</name></connection>
<intersection>271 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>265.5,14.5,265.5,15</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269.5,7.5,269.5,24.5</points>
<connection>
<GID>306</GID>
<name>OUT_0</name></connection>
<intersection>7.5 5</intersection>
<intersection>15 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>267.5,15,269.5,15</points>
<connection>
<GID>307</GID>
<name>IN_1</name></connection>
<intersection>269.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>269.5,7.5,271,7.5</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>269.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>458</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,9.5,270.5,26.5</points>
<intersection>9.5 1</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270.5,9.5,271,9.5</points>
<connection>
<GID>275</GID>
<name>IN_2</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>269.5,26.5,270.5,26.5</points>
<connection>
<GID>306</GID>
<name>OUT_2</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>459</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,8.5,270,25.5</points>
<intersection>8.5 3</intersection>
<intersection>25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>269.5,25.5,270,25.5</points>
<connection>
<GID>306</GID>
<name>OUT_1</name></connection>
<intersection>270 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>270,8.5,271,8.5</points>
<connection>
<GID>275</GID>
<name>IN_1</name></connection>
<intersection>270 0</intersection></hsegment></shape></wire>
<wire>
<ID>460</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,21,261,31</points>
<intersection>21 4</intersection>
<intersection>31 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>261,31,265.5,31</points>
<intersection>261 0</intersection>
<intersection>265.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>261,21,277,21</points>
<intersection>261 0</intersection>
<intersection>264.5 7</intersection>
<intersection>277 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>277,21,277,21.5</points>
<connection>
<GID>274</GID>
<name>OUT</name></connection>
<connection>
<GID>273</GID>
<name>clear</name></connection>
<intersection>21 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>264.5,21,264.5,21.5</points>
<connection>
<GID>306</GID>
<name>clock</name></connection>
<intersection>21 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>265.5,30.5,265.5,31</points>
<connection>
<GID>306</GID>
<name>count_enable</name></connection>
<intersection>31 3</intersection></vsegment></shape></wire>
<wire>
<ID>461</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,10.5,260.5,27.5</points>
<connection>
<GID>308</GID>
<name>IN_3</name></connection>
<intersection>14.5 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255,14.5,260.5,14.5</points>
<intersection>255 17</intersection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259,27.5,260.5,27.5</points>
<connection>
<GID>309</GID>
<name>OUT_3</name></connection>
<intersection>260.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>255,14.5,255,15</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>462</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259,7.5,259,24.5</points>
<connection>
<GID>309</GID>
<name>OUT_0</name></connection>
<intersection>7.5 5</intersection>
<intersection>15 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>257,15,259,15</points>
<connection>
<GID>310</GID>
<name>IN_1</name></connection>
<intersection>259 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>259,7.5,260.5,7.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>259 0</intersection></hsegment></shape></wire>
<wire>
<ID>463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,9.5,260,26.5</points>
<intersection>9.5 1</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,9.5,260.5,9.5</points>
<connection>
<GID>308</GID>
<name>IN_2</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259,26.5,260,26.5</points>
<connection>
<GID>309</GID>
<name>OUT_2</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>464</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,8.5,259.5,25.5</points>
<intersection>8.5 3</intersection>
<intersection>25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>259,25.5,259.5,25.5</points>
<connection>
<GID>309</GID>
<name>OUT_1</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>259.5,8.5,260.5,8.5</points>
<connection>
<GID>308</GID>
<name>IN_1</name></connection>
<intersection>259.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>465</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,21.5,250.5,31</points>
<intersection>21.5 4</intersection>
<intersection>31 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>250.5,31,255,31</points>
<intersection>250.5 0</intersection>
<intersection>255 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>250.5,21.5,266.5,21.5</points>
<connection>
<GID>309</GID>
<name>clock</name></connection>
<intersection>250.5 0</intersection>
<intersection>266.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>266.5,21,266.5,21.5</points>
<connection>
<GID>307</GID>
<name>OUT</name></connection>
<connection>
<GID>306</GID>
<name>clear</name></connection>
<intersection>21.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>255,30.5,255,31</points>
<connection>
<GID>309</GID>
<name>count_enable</name></connection>
<intersection>31 3</intersection></vsegment></shape></wire>
<wire>
<ID>467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,10.5,250,27.5</points>
<connection>
<GID>311</GID>
<name>IN_3</name></connection>
<intersection>14.5 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244.5,14.5,250,14.5</points>
<intersection>244.5 17</intersection>
<intersection>250 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>248.5,27.5,250,27.5</points>
<connection>
<GID>312</GID>
<name>OUT_3</name></connection>
<intersection>250 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>244.5,14.5,244.5,15</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>468</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,37,302.5,54</points>
<connection>
<GID>276</GID>
<name>IN_3</name></connection>
<intersection>41 1</intersection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>297,41,302.5,41</points>
<intersection>297 17</intersection>
<intersection>302.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301,54,302.5,54</points>
<connection>
<GID>277</GID>
<name>OUT_3</name></connection>
<intersection>302.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>297,41,297,41.5</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>41 1</intersection></vsegment></shape></wire>
<wire>
<ID>469</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301,34,301,51</points>
<connection>
<GID>277</GID>
<name>OUT_0</name></connection>
<intersection>34 5</intersection>
<intersection>41.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>299,41.5,301,41.5</points>
<connection>
<GID>278</GID>
<name>IN_1</name></connection>
<intersection>301 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>301,34,302.5,34</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>301 0</intersection></hsegment></shape></wire>
<wire>
<ID>470</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,36,302,53</points>
<intersection>36 1</intersection>
<intersection>53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302,36,302.5,36</points>
<connection>
<GID>276</GID>
<name>IN_2</name></connection>
<intersection>302 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301,53,302,53</points>
<connection>
<GID>277</GID>
<name>OUT_2</name></connection>
<intersection>302 0</intersection></hsegment></shape></wire>
<wire>
<ID>471</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,35,301.5,52</points>
<intersection>35 3</intersection>
<intersection>52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>301,52,301.5,52</points>
<connection>
<GID>277</GID>
<name>OUT_1</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>301.5,35,302.5,35</points>
<connection>
<GID>276</GID>
<name>IN_1</name></connection>
<intersection>301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>472</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298,47.5,298,48</points>
<connection>
<GID>278</GID>
<name>OUT</name></connection>
<connection>
<GID>277</GID>
<name>clear</name></connection>
<intersection>47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282,47.5,298,47.5</points>
<intersection>282 2</intersection>
<intersection>285.5 7</intersection>
<intersection>298 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>282,47.5,282,57.5</points>
<intersection>47.5 1</intersection>
<intersection>57.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>282,57.5,286.5,57.5</points>
<intersection>282 2</intersection>
<intersection>286.5 10</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>285.5,47.5,285.5,48</points>
<connection>
<GID>280</GID>
<name>clock</name></connection>
<intersection>47.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>286.5,57,286.5,57.5</points>
<connection>
<GID>280</GID>
<name>count_enable</name></connection>
<intersection>57.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>473</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248.5,7.5,248.5,24.5</points>
<connection>
<GID>312</GID>
<name>OUT_0</name></connection>
<intersection>7.5 5</intersection>
<intersection>15 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>246.5,15,248.5,15</points>
<connection>
<GID>313</GID>
<name>IN_1</name></connection>
<intersection>248.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>248.5,7.5,250,7.5</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>248.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>474</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,37,292,54</points>
<connection>
<GID>279</GID>
<name>IN_3</name></connection>
<intersection>41 1</intersection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286.5,41,292,41</points>
<intersection>286.5 17</intersection>
<intersection>292 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>290.5,54,292,54</points>
<connection>
<GID>280</GID>
<name>OUT_3</name></connection>
<intersection>292 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>286.5,41,286.5,41.5</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>41 1</intersection></vsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,34,290.5,51</points>
<connection>
<GID>280</GID>
<name>OUT_0</name></connection>
<intersection>34 5</intersection>
<intersection>41.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>288.5,41.5,290.5,41.5</points>
<connection>
<GID>281</GID>
<name>IN_1</name></connection>
<intersection>290.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>290.5,34,292,34</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>290.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,36,291.5,53</points>
<intersection>36 1</intersection>
<intersection>53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>291.5,36,292,36</points>
<connection>
<GID>279</GID>
<name>IN_2</name></connection>
<intersection>291.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>290.5,53,291.5,53</points>
<connection>
<GID>280</GID>
<name>OUT_2</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,35,291,52</points>
<intersection>35 3</intersection>
<intersection>52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>290.5,52,291,52</points>
<connection>
<GID>280</GID>
<name>OUT_1</name></connection>
<intersection>291 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>291,35,292,35</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<intersection>291 0</intersection></hsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287.5,47.5,287.5,48</points>
<connection>
<GID>281</GID>
<name>OUT</name></connection>
<connection>
<GID>280</GID>
<name>clear</name></connection>
<intersection>48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>271.5,48,287.5,48</points>
<connection>
<GID>283</GID>
<name>clock</name></connection>
<intersection>271.5 2</intersection>
<intersection>287.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>271.5,48,271.5,57.5</points>
<intersection>48 1</intersection>
<intersection>57.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>271.5,57.5,276,57.5</points>
<intersection>271.5 2</intersection>
<intersection>276 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>276,57,276,57.5</points>
<connection>
<GID>283</GID>
<name>count_enable</name></connection>
<intersection>57.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,37,281.5,54</points>
<connection>
<GID>282</GID>
<name>IN_3</name></connection>
<intersection>41 1</intersection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,41,281.5,41</points>
<intersection>276 17</intersection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280,54,281.5,54</points>
<connection>
<GID>283</GID>
<name>OUT_3</name></connection>
<intersection>281.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>276,41,276,41.5</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>41 1</intersection></vsegment></shape></wire>
<wire>
<ID>480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280,34,280,51</points>
<connection>
<GID>283</GID>
<name>OUT_0</name></connection>
<intersection>34 5</intersection>
<intersection>41.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>278,41.5,280,41.5</points>
<connection>
<GID>284</GID>
<name>IN_1</name></connection>
<intersection>280 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>280,34,281.5,34</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>280 0</intersection></hsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,36,281,53</points>
<intersection>36 1</intersection>
<intersection>53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281,36,281.5,36</points>
<connection>
<GID>282</GID>
<name>IN_2</name></connection>
<intersection>281 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280,53,281,53</points>
<connection>
<GID>283</GID>
<name>OUT_2</name></connection>
<intersection>281 0</intersection></hsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280.5,35,280.5,52</points>
<intersection>35 3</intersection>
<intersection>52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>280,52,280.5,52</points>
<connection>
<GID>283</GID>
<name>OUT_1</name></connection>
<intersection>280.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>280.5,35,281.5,35</points>
<connection>
<GID>282</GID>
<name>IN_1</name></connection>
<intersection>280.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,37,271,54</points>
<connection>
<GID>285</GID>
<name>IN_3</name></connection>
<intersection>41 1</intersection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>265.5,41,271,41</points>
<intersection>265.5 17</intersection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>269.5,54,271,54</points>
<connection>
<GID>286</GID>
<name>OUT_3</name></connection>
<intersection>271 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>265.5,41,265.5,41.5</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>41 1</intersection></vsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269.5,34,269.5,51</points>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection>
<intersection>34 5</intersection>
<intersection>41.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>267.5,41.5,269.5,41.5</points>
<connection>
<GID>287</GID>
<name>IN_1</name></connection>
<intersection>269.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>269.5,34,271,34</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>269.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,36,270.5,53</points>
<intersection>36 1</intersection>
<intersection>53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270.5,36,271,36</points>
<connection>
<GID>285</GID>
<name>IN_2</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>269.5,53,270.5,53</points>
<connection>
<GID>286</GID>
<name>OUT_2</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,35,270,52</points>
<intersection>35 3</intersection>
<intersection>52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>269.5,52,270,52</points>
<connection>
<GID>286</GID>
<name>OUT_1</name></connection>
<intersection>270 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>270,35,271,35</points>
<connection>
<GID>285</GID>
<name>IN_1</name></connection>
<intersection>270 0</intersection></hsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,47.5,261,57.5</points>
<intersection>47.5 4</intersection>
<intersection>57.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>261,57.5,265.5,57.5</points>
<intersection>261 0</intersection>
<intersection>265.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>261,47.5,277,47.5</points>
<intersection>261 0</intersection>
<intersection>264.5 7</intersection>
<intersection>277 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>277,47.5,277,48</points>
<connection>
<GID>284</GID>
<name>OUT</name></connection>
<connection>
<GID>283</GID>
<name>clear</name></connection>
<intersection>47.5 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>264.5,47.5,264.5,48</points>
<connection>
<GID>286</GID>
<name>clock</name></connection>
<intersection>47.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>265.5,57,265.5,57.5</points>
<connection>
<GID>286</GID>
<name>count_enable</name></connection>
<intersection>57.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,37,260.5,54</points>
<connection>
<GID>288</GID>
<name>IN_3</name></connection>
<intersection>41 1</intersection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255,41,260.5,41</points>
<intersection>255 17</intersection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259,54,260.5,54</points>
<connection>
<GID>289</GID>
<name>OUT_3</name></connection>
<intersection>260.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>255,41,255,41.5</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>41 1</intersection></vsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259,34,259,51</points>
<connection>
<GID>289</GID>
<name>OUT_0</name></connection>
<intersection>34 5</intersection>
<intersection>41.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>257,41.5,259,41.5</points>
<connection>
<GID>290</GID>
<name>IN_1</name></connection>
<intersection>259 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>259,34,260.5,34</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>259 0</intersection></hsegment></shape></wire>
<wire>
<ID>490</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,36,260,53</points>
<intersection>36 1</intersection>
<intersection>53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,36,260.5,36</points>
<connection>
<GID>288</GID>
<name>IN_2</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259,53,260,53</points>
<connection>
<GID>289</GID>
<name>OUT_2</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,35,259.5,52</points>
<intersection>35 3</intersection>
<intersection>52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>259,52,259.5,52</points>
<connection>
<GID>289</GID>
<name>OUT_1</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>259.5,35,260.5,35</points>
<connection>
<GID>288</GID>
<name>IN_1</name></connection>
<intersection>259.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,9.5,249.5,26.5</points>
<intersection>9.5 1</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>249.5,9.5,250,9.5</points>
<connection>
<GID>311</GID>
<name>IN_2</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>248.5,26.5,249.5,26.5</points>
<connection>
<GID>312</GID>
<name>OUT_2</name></connection>
<intersection>249.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,48,250.5,57.5</points>
<intersection>48 4</intersection>
<intersection>57.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>250.5,57.5,255,57.5</points>
<intersection>250.5 0</intersection>
<intersection>255 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>250.5,48,266.5,48</points>
<connection>
<GID>289</GID>
<name>clock</name></connection>
<intersection>250.5 0</intersection>
<intersection>266.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>266.5,47.5,266.5,48</points>
<connection>
<GID>287</GID>
<name>OUT</name></connection>
<connection>
<GID>286</GID>
<name>clear</name></connection>
<intersection>48 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>255,57,255,57.5</points>
<connection>
<GID>289</GID>
<name>count_enable</name></connection>
<intersection>57.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,48,292.5,57.5</points>
<intersection>48 4</intersection>
<intersection>57.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>292.5,57.5,297,57.5</points>
<intersection>292.5 0</intersection>
<intersection>297 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>292.5,48,296,48</points>
<connection>
<GID>277</GID>
<name>clock</name></connection>
<intersection>292.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>297,57,297,58.5</points>
<connection>
<GID>277</GID>
<name>count_enable</name></connection>
<intersection>57.5 3</intersection>
<intersection>58.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>196,58.5,297,58.5</points>
<intersection>196 7</intersection>
<intersection>297 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>196,21,196,58.5</points>
<intersection>21 8</intersection>
<intersection>58.5 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>196,21,203.5,21</points>
<connection>
<GID>325</GID>
<name>OUT</name></connection>
<intersection>196 7</intersection>
<intersection>203.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>203.5,21,203.5,21.5</points>
<connection>
<GID>324</GID>
<name>clear</name></connection>
<intersection>21 8</intersection></vsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,37,250,54</points>
<connection>
<GID>291</GID>
<name>IN_3</name></connection>
<intersection>41 1</intersection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244.5,41,250,41</points>
<intersection>244.5 17</intersection>
<intersection>250 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>248.5,54,250,54</points>
<connection>
<GID>292</GID>
<name>OUT_3</name></connection>
<intersection>250 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>244.5,41,244.5,41.5</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>41 1</intersection></vsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248.5,34,248.5,51</points>
<connection>
<GID>292</GID>
<name>OUT_0</name></connection>
<intersection>34 5</intersection>
<intersection>41.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>246.5,41.5,248.5,41.5</points>
<connection>
<GID>293</GID>
<name>IN_1</name></connection>
<intersection>248.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>248.5,34,250,34</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>248.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,36,249.5,53</points>
<intersection>36 1</intersection>
<intersection>53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>249.5,36,250,36</points>
<connection>
<GID>291</GID>
<name>IN_2</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>248.5,53,249.5,53</points>
<connection>
<GID>292</GID>
<name>OUT_2</name></connection>
<intersection>249.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249,35,249,52</points>
<intersection>35 3</intersection>
<intersection>52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>248.5,52,249,52</points>
<connection>
<GID>292</GID>
<name>OUT_1</name></connection>
<intersection>249 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>249,35,250,35</points>
<connection>
<GID>291</GID>
<name>IN_1</name></connection>
<intersection>249 0</intersection></hsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249,8.5,249,25.5</points>
<intersection>8.5 3</intersection>
<intersection>25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>248.5,25.5,249,25.5</points>
<connection>
<GID>312</GID>
<name>OUT_1</name></connection>
<intersection>249 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>249,8.5,250,8.5</points>
<connection>
<GID>311</GID>
<name>IN_1</name></connection>
<intersection>249 0</intersection></hsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239.5,37,239.5,54</points>
<connection>
<GID>294</GID>
<name>IN_3</name></connection>
<intersection>41 1</intersection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234,41,239.5,41</points>
<intersection>234 17</intersection>
<intersection>239.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238,54,239.5,54</points>
<connection>
<GID>295</GID>
<name>OUT_3</name></connection>
<intersection>239.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>234,41,234,41.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>41 1</intersection></vsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238,34,238,51</points>
<connection>
<GID>295</GID>
<name>OUT_0</name></connection>
<intersection>34 5</intersection>
<intersection>41.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>236,41.5,238,41.5</points>
<connection>
<GID>296</GID>
<name>IN_1</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>238,34,239.5,34</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>238 0</intersection></hsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,36,239,53</points>
<intersection>36 1</intersection>
<intersection>53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239,36,239.5,36</points>
<connection>
<GID>294</GID>
<name>IN_2</name></connection>
<intersection>239 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238,53,239,53</points>
<connection>
<GID>295</GID>
<name>OUT_2</name></connection>
<intersection>239 0</intersection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,35,238.5,52</points>
<intersection>35 3</intersection>
<intersection>52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>238,52,238.5,52</points>
<connection>
<GID>295</GID>
<name>OUT_1</name></connection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>238.5,35,239.5,35</points>
<connection>
<GID>294</GID>
<name>IN_1</name></connection>
<intersection>238.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,47.5,235,48</points>
<connection>
<GID>296</GID>
<name>OUT</name></connection>
<connection>
<GID>295</GID>
<name>clear</name></connection>
<intersection>47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,47.5,235,47.5</points>
<intersection>219 2</intersection>
<intersection>222.5 10</intersection>
<intersection>235 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>219,47.5,219,57.5</points>
<intersection>47.5 1</intersection>
<intersection>57.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>219,57.5,223.5,57.5</points>
<intersection>219 2</intersection>
<intersection>223.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>223.5,57,223.5,57.5</points>
<connection>
<GID>298</GID>
<name>count_enable</name></connection>
<intersection>57.5 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>222.5,47.5,222.5,48</points>
<connection>
<GID>298</GID>
<name>clock</name></connection>
<intersection>47.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,37,229,54</points>
<connection>
<GID>297</GID>
<name>IN_3</name></connection>
<intersection>41 1</intersection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>223.5,41,229,41</points>
<intersection>223.5 17</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227.5,54,229,54</points>
<connection>
<GID>298</GID>
<name>OUT_3</name></connection>
<intersection>229 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>223.5,41,223.5,41.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>41 1</intersection></vsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227.5,34,227.5,51</points>
<connection>
<GID>298</GID>
<name>OUT_0</name></connection>
<intersection>34 5</intersection>
<intersection>41.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>225.5,41.5,227.5,41.5</points>
<connection>
<GID>299</GID>
<name>IN_1</name></connection>
<intersection>227.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>227.5,34,229,34</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>227.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,36,228.5,53</points>
<intersection>36 1</intersection>
<intersection>53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>228.5,36,229,36</points>
<connection>
<GID>297</GID>
<name>IN_2</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227.5,53,228.5,53</points>
<connection>
<GID>298</GID>
<name>OUT_2</name></connection>
<intersection>228.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,35,228,52</points>
<intersection>35 3</intersection>
<intersection>52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>227.5,52,228,52</points>
<connection>
<GID>298</GID>
<name>OUT_1</name></connection>
<intersection>228 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>228,35,229,35</points>
<connection>
<GID>297</GID>
<name>IN_1</name></connection>
<intersection>228 0</intersection></hsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,37,218.5,54</points>
<connection>
<GID>300</GID>
<name>IN_3</name></connection>
<intersection>41 1</intersection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213,41,218.5,41</points>
<intersection>213 17</intersection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>217,54,218.5,54</points>
<connection>
<GID>301</GID>
<name>OUT_3</name></connection>
<intersection>218.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>213,41,213,41.5</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>41 1</intersection></vsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217,34,217,51</points>
<connection>
<GID>301</GID>
<name>OUT_0</name></connection>
<intersection>34 5</intersection>
<intersection>41.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>215,41.5,217,41.5</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>217,34,218.5,34</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,36,218,53</points>
<intersection>36 1</intersection>
<intersection>53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,36,218.5,36</points>
<connection>
<GID>300</GID>
<name>IN_2</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>217,53,218,53</points>
<connection>
<GID>301</GID>
<name>OUT_2</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217.5,35,217.5,52</points>
<intersection>35 3</intersection>
<intersection>52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>217,52,217.5,52</points>
<connection>
<GID>301</GID>
<name>OUT_1</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>217.5,35,218.5,35</points>
<connection>
<GID>300</GID>
<name>IN_1</name></connection>
<intersection>217.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>513</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,48,208.5,57.5</points>
<intersection>48 4</intersection>
<intersection>57.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>208.5,57.5,213,57.5</points>
<intersection>208.5 0</intersection>
<intersection>213 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>208.5,48,224.5,48</points>
<connection>
<GID>301</GID>
<name>clock</name></connection>
<intersection>208.5 0</intersection>
<intersection>224.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>224.5,47.5,224.5,48</points>
<connection>
<GID>299</GID>
<name>OUT</name></connection>
<connection>
<GID>298</GID>
<name>clear</name></connection>
<intersection>48 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>213,57,213,57.5</points>
<connection>
<GID>301</GID>
<name>count_enable</name></connection>
<intersection>57.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>514</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,37,208,54</points>
<connection>
<GID>303</GID>
<name>IN_3</name></connection>
<intersection>41 1</intersection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,41,208,41</points>
<intersection>202.5 17</intersection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>206.5,54,208,54</points>
<connection>
<GID>304</GID>
<name>OUT_3</name></connection>
<intersection>208 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>202.5,41,202.5,41.5</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>41 1</intersection></vsegment></shape></wire>
<wire>
<ID>515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,34,206.5,51</points>
<connection>
<GID>304</GID>
<name>OUT_0</name></connection>
<intersection>34 5</intersection>
<intersection>41.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>204.5,41.5,206.5,41.5</points>
<connection>
<GID>305</GID>
<name>IN_1</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>206.5,34,208,34</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>206.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,36,207.5,53</points>
<intersection>36 1</intersection>
<intersection>53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207.5,36,208,36</points>
<connection>
<GID>303</GID>
<name>IN_2</name></connection>
<intersection>207.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>206.5,53,207.5,53</points>
<connection>
<GID>304</GID>
<name>OUT_2</name></connection>
<intersection>207.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,35,207,52</points>
<intersection>35 3</intersection>
<intersection>52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>206.5,52,207,52</points>
<connection>
<GID>304</GID>
<name>OUT_1</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>207,35,208,35</points>
<connection>
<GID>303</GID>
<name>IN_1</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203.5,47.5,203.5,48</points>
<connection>
<GID>305</GID>
<name>OUT</name></connection>
<connection>
<GID>304</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>519</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198,47.5,198,57.5</points>
<intersection>47.5 4</intersection>
<intersection>57.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,57.5,202.5,57.5</points>
<intersection>198 0</intersection>
<intersection>202.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>198,47.5,214,47.5</points>
<intersection>198 0</intersection>
<intersection>201.5 15</intersection>
<intersection>214 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>214,47.5,214,48</points>
<connection>
<GID>302</GID>
<name>OUT</name></connection>
<connection>
<GID>301</GID>
<name>clear</name></connection>
<intersection>47.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>202.5,57,202.5,57.5</points>
<connection>
<GID>304</GID>
<name>count_enable</name></connection>
<intersection>57.5 3</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>201.5,47.5,201.5,48</points>
<connection>
<GID>304</GID>
<name>clock</name></connection>
<intersection>47.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239.5,10.5,239.5,27.5</points>
<connection>
<GID>314</GID>
<name>IN_3</name></connection>
<intersection>14.5 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234,14.5,239.5,14.5</points>
<intersection>234 17</intersection>
<intersection>239.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238,27.5,239.5,27.5</points>
<connection>
<GID>315</GID>
<name>OUT_3</name></connection>
<intersection>239.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>234,14.5,234,15</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>256,47.5,256,48</points>
<connection>
<GID>290</GID>
<name>OUT</name></connection>
<connection>
<GID>289</GID>
<name>clear</name></connection>
<intersection>47.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>240,47.5,256,47.5</points>
<intersection>240 4</intersection>
<intersection>243.5 8</intersection>
<intersection>256 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>240,47.5,240,57.5</points>
<intersection>47.5 3</intersection>
<intersection>57.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>240,57.5,244.5,57.5</points>
<intersection>240 4</intersection>
<intersection>244.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>244.5,57,244.5,57.5</points>
<connection>
<GID>292</GID>
<name>count_enable</name></connection>
<intersection>57.5 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>243.5,47.5,243.5,48</points>
<connection>
<GID>292</GID>
<name>clock</name></connection>
<intersection>47.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,47.5,245.5,48</points>
<connection>
<GID>293</GID>
<name>OUT</name></connection>
<connection>
<GID>292</GID>
<name>clear</name></connection>
<intersection>48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229.5,48,245.5,48</points>
<connection>
<GID>295</GID>
<name>clock</name></connection>
<intersection>229.5 4</intersection>
<intersection>245.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>229.5,48,229.5,57.5</points>
<intersection>48 1</intersection>
<intersection>57.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>229.5,57.5,234,57.5</points>
<intersection>229.5 4</intersection>
<intersection>234 17</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>234,57,234,57.5</points>
<connection>
<GID>295</GID>
<name>count_enable</name></connection>
<intersection>57.5 15</intersection></vsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238,7.5,238,24.5</points>
<connection>
<GID>315</GID>
<name>OUT_0</name></connection>
<intersection>7.5 5</intersection>
<intersection>15 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>236,15,238,15</points>
<connection>
<GID>316</GID>
<name>IN_1</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>238,7.5,239.5,7.5</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>238 0</intersection></hsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,9.5,239,26.5</points>
<intersection>9.5 1</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239,9.5,239.5,9.5</points>
<connection>
<GID>314</GID>
<name>IN_2</name></connection>
<intersection>239 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238,26.5,239,26.5</points>
<connection>
<GID>315</GID>
<name>OUT_2</name></connection>
<intersection>239 0</intersection></hsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,8.5,238.5,25.5</points>
<intersection>8.5 3</intersection>
<intersection>25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>238,25.5,238.5,25.5</points>
<connection>
<GID>315</GID>
<name>OUT_1</name></connection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>238.5,8.5,239.5,8.5</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<intersection>238.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,21,235,21.5</points>
<connection>
<GID>316</GID>
<name>OUT</name></connection>
<connection>
<GID>315</GID>
<name>clear</name></connection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,21,235,21</points>
<intersection>219 2</intersection>
<intersection>222.5 10</intersection>
<intersection>235 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>219,21,219,31</points>
<intersection>21 1</intersection>
<intersection>31 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>219,31,223.5,31</points>
<intersection>219 2</intersection>
<intersection>223.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>223.5,30.5,223.5,31</points>
<connection>
<GID>318</GID>
<name>count_enable</name></connection>
<intersection>31 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>222.5,21,222.5,21.5</points>
<connection>
<GID>318</GID>
<name>clock</name></connection>
<intersection>21 1</intersection></vsegment></shape></wire>
<wire>
<ID>527</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,10.5,229,27.5</points>
<connection>
<GID>317</GID>
<name>IN_3</name></connection>
<intersection>14.5 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>223.5,14.5,229,14.5</points>
<intersection>223.5 17</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227.5,27.5,229,27.5</points>
<connection>
<GID>318</GID>
<name>OUT_3</name></connection>
<intersection>229 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>223.5,14.5,223.5,15</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>528</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227.5,7.5,227.5,24.5</points>
<connection>
<GID>318</GID>
<name>OUT_0</name></connection>
<intersection>7.5 5</intersection>
<intersection>15 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>225.5,15,227.5,15</points>
<connection>
<GID>319</GID>
<name>IN_1</name></connection>
<intersection>227.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>227.5,7.5,229,7.5</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>227.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,9.5,228.5,26.5</points>
<intersection>9.5 1</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>228.5,9.5,229,9.5</points>
<connection>
<GID>317</GID>
<name>IN_2</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227.5,26.5,228.5,26.5</points>
<connection>
<GID>318</GID>
<name>OUT_2</name></connection>
<intersection>228.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,8.5,228,25.5</points>
<intersection>8.5 3</intersection>
<intersection>25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>227.5,25.5,228,25.5</points>
<connection>
<GID>318</GID>
<name>OUT_1</name></connection>
<intersection>228 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>228,8.5,229,8.5</points>
<connection>
<GID>317</GID>
<name>IN_1</name></connection>
<intersection>228 0</intersection></hsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,10.5,218.5,27.5</points>
<connection>
<GID>320</GID>
<name>IN_3</name></connection>
<intersection>14.5 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213,14.5,218.5,14.5</points>
<intersection>213 17</intersection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>217,27.5,218.5,27.5</points>
<connection>
<GID>321</GID>
<name>OUT_3</name></connection>
<intersection>218.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>213,14.5,213,15</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217,7.5,217,24.5</points>
<connection>
<GID>321</GID>
<name>OUT_0</name></connection>
<intersection>7.5 5</intersection>
<intersection>15 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>215,15,217,15</points>
<connection>
<GID>322</GID>
<name>IN_1</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>217,7.5,218.5,7.5</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,9.5,218,26.5</points>
<intersection>9.5 1</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,9.5,218.5,9.5</points>
<connection>
<GID>320</GID>
<name>IN_2</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>217,26.5,218,26.5</points>
<connection>
<GID>321</GID>
<name>OUT_2</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>534</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217.5,8.5,217.5,25.5</points>
<intersection>8.5 3</intersection>
<intersection>25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>217,25.5,217.5,25.5</points>
<connection>
<GID>321</GID>
<name>OUT_1</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>217.5,8.5,218.5,8.5</points>
<connection>
<GID>320</GID>
<name>IN_1</name></connection>
<intersection>217.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>535</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,21.5,208.5,31</points>
<intersection>21.5 4</intersection>
<intersection>31 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>208.5,31,213,31</points>
<intersection>208.5 0</intersection>
<intersection>213 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>208.5,21.5,224.5,21.5</points>
<connection>
<GID>321</GID>
<name>clock</name></connection>
<intersection>208.5 0</intersection>
<intersection>224.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>224.5,21,224.5,21.5</points>
<connection>
<GID>319</GID>
<name>OUT</name></connection>
<connection>
<GID>318</GID>
<name>clear</name></connection>
<intersection>21.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>213,30.5,213,31</points>
<connection>
<GID>321</GID>
<name>count_enable</name></connection>
<intersection>31 3</intersection></vsegment></shape></wire>
<wire>
<ID>536</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,10.5,208,27.5</points>
<connection>
<GID>323</GID>
<name>IN_3</name></connection>
<intersection>14.5 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,14.5,208,14.5</points>
<intersection>202.5 17</intersection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>206.5,27.5,208,27.5</points>
<connection>
<GID>324</GID>
<name>OUT_3</name></connection>
<intersection>208 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>202.5,14.5,202.5,15</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>537</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,7.5,206.5,24.5</points>
<connection>
<GID>324</GID>
<name>OUT_0</name></connection>
<intersection>7.5 5</intersection>
<intersection>15 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>204.5,15,206.5,15</points>
<connection>
<GID>325</GID>
<name>IN_1</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>206.5,7.5,208,7.5</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>206.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>538</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,9.5,207.5,26.5</points>
<intersection>9.5 1</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207.5,9.5,208,9.5</points>
<connection>
<GID>323</GID>
<name>IN_2</name></connection>
<intersection>207.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>206.5,26.5,207.5,26.5</points>
<connection>
<GID>324</GID>
<name>OUT_2</name></connection>
<intersection>207.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>539</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,8.5,207,25.5</points>
<intersection>8.5 3</intersection>
<intersection>25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>206.5,25.5,207,25.5</points>
<connection>
<GID>324</GID>
<name>OUT_1</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>207,8.5,208,8.5</points>
<connection>
<GID>323</GID>
<name>IN_1</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>540</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198,21,198,31</points>
<intersection>21 4</intersection>
<intersection>31 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,31,202.5,31</points>
<intersection>198 0</intersection>
<intersection>202.5 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>198,21,214,21</points>
<intersection>198 0</intersection>
<intersection>201.5 15</intersection>
<intersection>214 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>214,21,214,21.5</points>
<connection>
<GID>322</GID>
<name>OUT</name></connection>
<connection>
<GID>321</GID>
<name>clear</name></connection>
<intersection>21 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>202.5,30.5,202.5,31</points>
<connection>
<GID>324</GID>
<name>count_enable</name></connection>
<intersection>31 3</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>201.5,21,201.5,21.5</points>
<connection>
<GID>324</GID>
<name>clock</name></connection>
<intersection>21 4</intersection></vsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>256,21,256,21.5</points>
<connection>
<GID>310</GID>
<name>OUT</name></connection>
<connection>
<GID>309</GID>
<name>clear</name></connection>
<intersection>21 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>240,21,256,21</points>
<intersection>240 4</intersection>
<intersection>243.5 8</intersection>
<intersection>256 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>240,21,240,31</points>
<intersection>21 3</intersection>
<intersection>31 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>240,31,244.5,31</points>
<intersection>240 4</intersection>
<intersection>244.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>244.5,30.5,244.5,31</points>
<connection>
<GID>312</GID>
<name>count_enable</name></connection>
<intersection>31 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>243.5,21,243.5,21.5</points>
<connection>
<GID>312</GID>
<name>clock</name></connection>
<intersection>21 3</intersection></vsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,21,245.5,21.5</points>
<connection>
<GID>313</GID>
<name>OUT</name></connection>
<connection>
<GID>312</GID>
<name>clear</name></connection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229.5,21,245.5,21</points>
<intersection>229.5 4</intersection>
<intersection>233 20</intersection>
<intersection>245.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>229.5,21,229.5,30.5</points>
<intersection>21 1</intersection>
<intersection>30.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>229.5,30.5,234,30.5</points>
<connection>
<GID>315</GID>
<name>count_enable</name></connection>
<intersection>229.5 4</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>233,21,233,21.5</points>
<connection>
<GID>315</GID>
<name>clock</name></connection>
<intersection>21 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-2.72885,92.3199,1406,-634.228</PageViewport></page 1>
<page 2>
<PageViewport>-2.72885,92.3199,1406,-634.228</PageViewport></page 2>
<page 3>
<PageViewport>-2.72885,92.3199,1406,-634.228</PageViewport></page 3>
<page 4>
<PageViewport>-2.72885,92.3199,1406,-634.228</PageViewport></page 4>
<page 5>
<PageViewport>-2.72885,92.3199,1406,-634.228</PageViewport></page 5>
<page 6>
<PageViewport>-2.72885,92.3199,1406,-634.228</PageViewport></page 6>
<page 7>
<PageViewport>-2.72885,92.3199,1406,-634.228</PageViewport></page 7>
<page 8>
<PageViewport>-2.72885,92.3199,1406,-634.228</PageViewport></page 8>
<page 9>
<PageViewport>-2.72885,92.3199,1406,-634.228</PageViewport></page 9></circuit>